MACRO gf180mcu_mux
    CLASS BLOCK BLACKBOX ;
    FOREIGN gf180mcu_mux ;
    ORIGIN 0.43 2.17 ;
    SIZE 17.37 BY 13.54 ;
    PIN z 
        PORT 
            LAYER Metal1 ;
                POLYGON 6.565 3.845 6.565 4.235 6.620 4.235 6.620 4.840 8.300 4.840 8.300 4.870 8.560 4.870 8.560 4.840 10.240 4.840 10.240 4.335 10.295 4.335 10.295 3.945 10.125 3.945 9.955 3.945 9.955 4.335 10.010 4.335 10.010 4.610 8.560 4.610 8.560 4.580 8.300 4.580 8.300 4.610 6.850 4.610 6.850 4.235 6.905 4.235 6.905 3.845 ;
                POLYGON 9.105 4.725 9.105 11.370 16.510 11.370 16.510 11.200 16.510 11.030 9.445 11.030 9.445 4.725 ;
        END 
    END z 
    PIN s0 
        PORT 
            LAYER Metal1 ;
                POLYGON 10.510 4.780 10.510 4.780 10.900 4.780 10.970 4.780 10.970 4.780 10.995 4.780 10.995 9.200 16.510 9.200 16.510 9.030 16.510 8.860 11.335 8.860 11.335 4.780 11.360 4.780 11.360 4.440 11.165 4.440 10.970 4.440 10.510 4.440 ;
        END 
    END s0 
    PIN s1b 
        PORT 
            LAYER Metal1 ;
                POLYGON 7.595 5.195 7.595 6.890 7.595 11.030 0 11.030 0 11.200 0 11.370 7.935 11.370 7.935 6.890 7.935 5.195 ;
        END 
    END s1b 
    PIN i1_r 
        PORT 
            LAYER Metal1 ;
                POLYGON 16.510 7.030 16.120 7.030 16.120 6.975 11.885 6.975 11.885 5.065 11.885 4.340 11.885 4.145 12.055 4.145 12.225 4.145 12.225 4.340 12.225 5.065 12.225 6.745 16.120 6.745 16.120 6.690 16.510 6.690 ;
        END 
    END i1_r 
    PIN i0_r 
        PORT 
            LAYER Metal1 ;
                POLYGON 14.285 3.650 14.285 4.090 14.285 4.460 14.115 4.460 16.120 4.460 16.510 4.460 16.510 4.630 16.510 4.800 16.510 4.800 16.315 4.800 13.945 4.800 13.945 4.090 13.945 3.650 ;
        END 
    END i0_r 
    PIN s1 
        PORT 
            LAYER Metal1 ;
                POLYGON 9.015 2.150 9.015 0.915 9.015 -2.170 0 -2.170 0 -2.000 0 -1.830 8.675 -1.830 8.675 0.915 8.675 2.150 ;
        END 
    END s1 
    PIN i3_r 
        PORT 
            LAYER Metal1 ;
                POLYGON 16.510 0.340 16.120 0.340 16.120 0.285 12.225 0.285 12.225 1.970 12.225 2.700 12.225 2.895 12.055 2.895 11.885 2.895 11.885 2.700 11.885 1.970 11.885 0.055 16.120 0.055 16.120 0 16.510 0 ;
        END 
    END i3_r 
    PIN i2_r 
        PORT 
            LAYER Metal1 ;
                POLYGON 13.945 3.390 13.945 2.945 13.945 2.230 14.115 2.230 16.120 2.230 16.510 2.230 16.510 2.400 16.510 2.570 16.510 2.570 16.315 2.570 14.285 2.570 14.285 2.945 14.285 3.390 ;
        END 
    END i2_r 
    PIN i1_l 
        PORT 
            LAYER Metal1 ;
                POLYGON 0 6.940 0.390 6.940 0.390 6.885 4.825 6.885 4.825 4.970 4.825 4.240 4.825 4.045 4.655 4.045 4.485 4.045 4.485 4.240 4.485 4.970 4.485 6.655 0.390 6.655 0.390 6.600 0 6.600 ;
        END 
    END i1_l 
    PIN s0b 
        PORT 
            LAYER Metal1 ;
                POLYGON 6.250 4.610 6.250 4.610 5.860 4.610 5.400 4.610 5.400 4.950 5.425 4.950 5.425 8.860 0 8.860 0 9.030 0 9.200 5.765 9.200 5.765 4.950 5.790 4.950 5.790 4.950 5.595 4.950 5.790 4.950 6.250 4.950 ;
        END 
    END s0b 
    PIN i3_l 
        PORT 
            LAYER Metal1 ;
                POLYGON 0 0.340 0.390 0.340 0.390 0.285 4.485 0.285 4.485 1.970 4.485 2.700 4.485 2.895 4.655 2.895 4.825 2.895 4.825 2.700 4.825 1.970 4.825 0.055 0.390 0.055 0.390 0 0 0 ;
        END 
    END i3_l 
    PIN i0_l 
        PORT 
            LAYER Metal1 ;
                POLYGON 2.225 3.950 2.225 4.300 2.225 4.400 2.395 4.400 0.390 4.400 0 4.400 0 4.570 0 4.740 0 4.740 0.195 4.740 2.565 4.740 2.565 4.300 2.565 3.950 ;
        END 
    END i0_l 
    PIN i2_l 
        PORT 
            LAYER Metal1 ;
                POLYGON 2.565 2.990 2.565 2.640 2.565 2.200 2.395 2.200 0.390 2.200 0 2.200 0 2.370 0 2.540 0 2.540 0.195 2.540 2.225 2.540 2.225 2.640 2.225 2.990 ;
        END 
    END i2_l 
    OBS 
        LAYER Metal1 ;
            POLYGON 3.330 4.315 3.330 4.315 4.255 4.315 4.255 3.815 5.055 3.815 5.055 4.160 5.170 4.160 5.410 4.160 5.800 4.160 5.800 3.990 5.800 3.820 5.800 3.820 5.605 3.820 5.285 3.820 5.285 3.585 4.025 3.585 4.025 3.975 4.140 3.975 3.330 3.975 ;
            POLYGON 3.355 2.600 3.355 2.955 3.355 3.355 7.695 3.355 7.695 3.705 7.695 3.995 7.695 4.190 7.865 4.190 8.035 4.190 8.035 3.995 8.035 3.705 8.035 3.125 3.695 3.125 3.695 2.955 3.695 2.600 ;
            POLYGON 13.280 4.015 13.280 4.015 12.455 4.015 12.455 3.915 11.655 3.915 11.655 4.060 11.540 4.060 11.350 4.060 10.960 4.060 10.960 3.890 10.960 3.720 10.960 3.720 11.155 3.720 11.425 3.720 11.425 3.685 12.685 3.685 12.685 3.675 12.570 3.675 13.280 3.675 ;
            POLYGON 13.255 3.000 13.255 3.390 12.915 3.390 12.915 3.355 9.265 3.355 9.265 3.630 9.265 3.895 9.265 4.090 9.095 4.090 8.925 4.090 8.925 3.895 8.925 3.630 8.925 3.125 12.915 3.125 12.915 3.090 12.915 3.090 12.915 3.000 ;
    END 
END gf180mcu_mux 
END LIBRARY 
