MACRO gf180mcu_mux ; 
    PIN s0 
        PORT 
            LAYER Metal1 ;
                POLYGON 8.510 2.780 8.510 2.780 8.625 2.780 9.015 2.780 9.015 2.610 9.015 2.440 9.015 2.440 8.900 2.440 8.510 2.440 ;
        END 
    END s0 
    PIN s0b 
        PORT 
            LAYER Metal1 ;
                POLYGON 4.250 2.610 4.250 2.610 4.135 2.610 3.745 2.610 3.745 2.780 3.745 2.950 3.745 2.950 3.860 2.950 4.250 2.950 ;
        END 
    END s0b 
    PIN i1 
        PORT 
            LAYER Metal1 ;
                POLYGON 0 2.938 0.390 2.938 0.390 2.883 2.825 2.883 2.825 2.469 2.825 2.240 2.825 2.045 2.655 2.045 2.485 2.045 2.485 2.240 2.485 2.469 2.485 2.653 0.390 2.653 0.390 2.598 0 2.598 ;
                POLYGON 12.510 3.040 12.120 3.040 12.120 2.985 9.885 2.985 9.885 2.570 9.885 2.340 9.885 2.145 10.055 2.145 10.225 2.145 10.225 2.340 10.225 2.570 10.225 2.755 12.120 2.755 12.120 2.700 12.510 2.700 ;
        END 
    END i1 
    PIN i0 
        PORT 
            LAYER Metal1 ;
                POLYGON 0.565 2.340 0.565 1.950 0.510 1.950 0.510 1.787 0.390 1.787 0.390 1.732 0 1.732 0 1.902 0 2.072 0.390 2.072 0.390 2.017 0.280 2.017 0.280 1.950 0.225 1.950 0.225 2.340 ;
                POLYGON 12.285 1.650 12.285 1.800 12.115 1.800 12.510 1.800 12.510 1.970 12.510 2.140 12.510 2.140 11.945 2.140 11.945 1.650 ;
        END 
    END i0 
    PIN i3 
        PORT 
            LAYER Metal1 ;
                POLYGON 0 0.340 0.390 0.340 0.390 0.285 2.485 0.285 2.485 0.470 2.485 0.700 2.485 0.895 2.655 0.895 2.825 0.895 2.825 0.700 2.825 0.470 2.825 0.055 0.390 0.055 0.390 0 0 0 ;
                POLYGON 12.510 0.340 12.120 0.340 12.120 0.285 10.225 0.285 10.225 0.470 10.225 0.700 10.225 0.895 10.055 0.895 9.885 0.895 9.885 0.700 9.885 0.470 9.885 0.055 12.120 0.055 12.120 0 12.510 0 ;
        END 
    END i3 
    PIN z 
        PORT 
            LAYER Metal1 ;
        END 
    END z 
    PIN i2 
        PORT 
            LAYER Metal1 ;
                POLYGON 0.225 0.600 0.225 0.990 0.280 0.990 0.280 0.921 0.390 0.921 0.390 0.866 0 0.866 0 1.036 0 1.206 0.390 1.206 0.390 1.151 0.510 1.151 0.510 0.990 0.565 0.990 0.565 0.600 ;
                POLYGON 11.945 1.390 11.945 0.900 12.115 0.900 12.510 0.900 12.510 1.070 12.510 1.240 12.510 1.240 12.285 1.240 12.285 1.390 ;
        END 
    END i2 
    PIN s1 
        PORT 
            LAYER Metal1 ;
                RECT 6.650 -0.240 7.040 0.150 ; 
        END 
    END s1 
    OBS 
        LAYER Metal1 ;
            POLYGON 1.330 2.315 1.330 2.315 2.255 2.315 2.255 1.815 3.055 1.815 3.055 2.162 3.170 2.162 3.410 2.162 3.800 2.162 3.800 1.992 3.800 1.822 3.800 1.822 3.605 1.822 3.285 1.822 3.285 1.585 2.025 1.585 2.025 1.975 2.140 1.975 1.330 1.975 ;
            POLYGON 1.355 0.600 1.355 0.955 1.355 1.355 5.695 1.355 5.695 1.707 5.695 1.993 5.695 2.188 5.865 2.188 6.035 2.188 6.035 1.993 6.035 1.707 6.035 1.125 1.695 1.125 1.695 0.955 1.695 0.600 ;
            POLYGON 11.280 2.015 11.280 2.015 10.455 2.015 10.455 1.915 9.655 1.915 9.655 2.062 9.540 2.062 9.350 2.062 8.960 2.062 8.960 1.892 8.960 1.722 8.960 1.722 9.155 1.722 9.425 1.722 9.425 1.685 10.685 1.685 10.685 1.675 10.570 1.675 11.280 1.675 ;
            POLYGON 11.255 1.000 11.255 1.390 10.915 1.390 10.915 1.355 7.265 1.355 7.265 1.632 7.265 1.893 7.265 2.088 7.095 2.088 6.925 2.088 6.925 1.893 6.925 1.632 6.925 1.125 10.915 1.125 10.915 1.090 10.915 1.090 10.915 1.000 ;
            POLYGON 4.565 1.845 4.565 2.235 4.620 2.235 4.620 2.842 6.300 2.842 6.300 2.872 6.560 2.872 6.560 2.842 8.240 2.842 8.240 2.335 8.295 2.335 8.295 1.945 8.125 1.945 7.955 1.945 7.955 2.335 8.010 2.335 8.010 2.612 6.560 2.612 6.560 2.582 6.300 2.582 6.300 2.612 4.850 2.612 4.850 2.235 4.905 2.235 4.905 1.845 ;
    END 
END gf180mcu_mux 
END LIBRARY 

