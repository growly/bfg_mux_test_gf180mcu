MACRO gf180mcu_mux
    CLASS BLOCK BLACKBOX ;
    FOREIGN gf180mcu_mux ;
    ORIGIN 0.45 0.31 ;
    SIZE 13.49 BY 3.92 ;
    PIN s0 
        PORT 
            LAYER Metal1 ;
                POLYGON 8.440 2.760 8.440 2.760 8.820 2.760 9.100 2.760 9.480 2.760 9.480 2.595 9.480 2.430 9.480 2.430 9.290 2.430 9.100 2.430 8.440 2.430 ;
        END 
    END s0 
    PIN z 
        PORT 
            LAYER Metal1 ;
                POLYGON 4.525 1.825 4.525 2.205 4.575 2.205 4.575 2.800 6.245 2.800 6.245 2.825 6.495 2.825 6.495 2.800 8.165 2.800 8.165 2.325 8.215 2.325 8.215 1.945 8.050 1.945 7.885 1.945 7.885 2.325 7.935 2.325 7.935 2.570 6.495 2.570 6.495 2.545 6.245 2.545 6.245 2.570 4.805 2.570 4.805 2.205 4.855 2.205 4.855 1.825 ;
        END 
    END z 
    PIN i0_r 
        PORT 
            LAYER Metal1 ;
                POLYGON 12.165 1.640 12.165 1.790 12.000 1.790 12.045 1.790 12.390 1.790 12.390 1.955 12.390 2.120 12.390 2.120 12.200 2.120 11.835 2.120 11.835 1.640 ;
        END 
    END i0_r 
    PIN i2_r 
        PORT 
            LAYER Metal1 ;
                POLYGON 11.835 1.380 11.835 0.895 12.000 0.895 12.045 0.895 12.390 0.895 12.390 1.060 12.390 1.225 12.390 1.225 12.200 1.225 12.165 1.225 12.165 1.380 ;
        END 
    END i2_r 
    PIN i1_l 
        PORT 
            LAYER Metal1 ;
                POLYGON 0 2.895 0.380 2.895 0.380 2.845 2.795 2.845 2.795 2.435 2.795 2.215 2.795 2.025 2.630 2.025 2.465 2.025 2.465 2.215 2.465 2.435 2.465 2.615 0.380 2.615 0.380 2.565 0 2.565 ;
        END 
    END i1_l 
    PIN s0b 
        PORT 
            LAYER Metal1 ;
                POLYGON 4.200 2.590 4.200 2.590 3.820 2.590 3.540 2.590 3.160 2.590 3.160 2.755 3.160 2.920 3.160 2.920 3.350 2.920 3.540 2.920 4.200 2.920 ;
        END 
    END s0b 
    PIN i3_l 
        PORT 
            LAYER Metal1 ;
                POLYGON 0 0.330 0.380 0.330 0.380 0.280 2.465 0.280 2.465 0.460 2.465 0.685 2.465 0.875 2.630 0.875 2.795 0.875 2.795 0.685 2.795 0.460 2.795 0.050 0.380 0.050 0.380 0 0 0 ;
        END 
    END i3_l 
    PIN i0_l 
        PORT 
            LAYER Metal1 ;
                POLYGON 0.555 2.300 0.555 2.000 0.555 1.710 0.390 1.710 0.380 1.710 0 1.710 0 1.875 0 2.040 0 2.040 0.190 2.040 0.225 2.040 0.225 2.000 0.225 2.300 ;
        END 
    END i0_l 
    PIN i2_l 
        PORT 
            LAYER Metal1 ;
                POLYGON 0.225 0.600 0.225 0.895 0.225 0.855 0.390 0.855 0.380 0.855 0 0.855 0 1.020 0 1.185 0 1.185 0.190 1.185 0.555 1.185 0.555 0.895 0.555 0.600 ;
        END 
    END i2_l 
    PIN i1_r 
        PORT 
            LAYER Metal1 ;
                POLYGON 12.390 3.015 12.010 3.015 12.010 2.965 9.795 2.965 9.795 2.555 9.795 2.335 9.795 2.145 9.960 2.145 10.125 2.145 10.125 2.335 10.125 2.555 10.125 2.735 12.010 2.735 12.010 2.685 12.390 2.685 ;
        END 
    END i1_r 
    PIN s1b 
        PORT 
            LAYER Metal1 ;
                RECT 5.520 3.165 5.900 3.545 ; 
        END 
    END s1b 
    PIN i3_r 
        PORT 
            LAYER Metal1 ;
                POLYGON 12.390 0.330 12.010 0.330 12.010 0.280 10.125 0.280 10.125 0.460 10.125 0.685 10.125 0.875 9.960 0.875 9.795 0.875 9.795 0.685 9.795 0.460 9.795 0.050 12.010 0.050 12.010 0 12.390 0 ;
        END 
    END i3_r 
    PIN s1 
        PORT 
            LAYER Metal1 ;
                RECT 6.590 -0.245 6.970 0.135 ; 
        END 
    END s1 
    OBS 
        LAYER Metal1 ;
            POLYGON 1.320 2.275 1.320 2.275 2.235 2.275 2.235 1.795 3.025 1.795 3.025 2.125 3.140 2.125 3.380 2.125 3.760 2.125 3.760 1.960 3.760 1.795 3.760 1.795 3.570 1.795 3.255 1.795 3.255 1.565 2.005 1.565 2.005 1.945 2.120 1.945 1.320 1.945 ;
            POLYGON 1.345 0.600 1.345 0.945 1.345 1.335 5.645 1.335 5.645 1.680 5.645 1.965 5.645 2.155 5.810 2.155 5.975 2.155 5.975 1.965 5.975 1.680 5.975 1.105 1.675 1.105 1.675 0.945 1.675 0.600 ;
            POLYGON 11.170 1.995 11.170 1.995 10.355 1.995 10.355 1.915 9.565 1.915 9.565 2.045 9.450 2.045 9.260 2.045 8.880 2.045 8.880 1.880 8.880 1.715 8.880 1.715 9.070 1.715 9.335 1.715 9.335 1.685 10.585 1.685 10.585 1.665 10.470 1.665 11.170 1.665 ;
            POLYGON 11.145 1.000 11.145 1.380 10.815 1.380 10.815 1.335 7.195 1.335 7.195 1.620 7.195 1.885 7.195 2.075 7.030 2.075 6.865 2.075 6.865 1.885 6.865 1.620 6.865 1.105 10.815 1.105 10.815 1.060 10.815 1.060 10.815 1.000 ;
    END 
END gf180mcu_mux 
END LIBRARY 
