(* blackbox *)
module gf180mcu_mux(
  input i0_l,
  input i1_l,
  input i2_l,
  input i3_l,
  input i0_r,
  input i1_r,
  input i2_r,
  input i3_r,
  input s0,
  input s0b,
  input s1,
  input s1b,
  output z
);
endmodule
