magic
tech gf180mcuC
magscale 1 5
timestamp 1670835587
<< obsm1 >>
rect 672 1538 14360 8262
<< metal2 >>
rect 2352 9600 2408 9900
rect 8736 9600 8792 9900
rect 14784 9600 14840 9900
rect 0 100 56 400
rect 6048 100 6104 400
rect 12432 100 12488 400
<< obsm2 >>
rect 14 9570 2322 9600
rect 2438 9570 8706 9600
rect 8822 9570 14754 9600
rect 14 430 14826 9570
rect 86 400 6018 430
rect 6134 400 12402 430
rect 12518 400 14826 430
<< metal3 >>
rect 100 6048 400 6104
rect 14600 3696 14900 3752
<< obsm3 >>
rect 9 6134 14831 8890
rect 9 6018 70 6134
rect 430 6018 14831 6134
rect 9 3782 14831 6018
rect 9 3666 14570 3782
rect 9 1246 14831 3666
<< metal4 >>
rect 2293 1538 2453 8262
rect 3994 1538 4154 8262
rect 5695 1538 5855 8262
rect 7396 1538 7556 8262
rect 9097 1538 9257 8262
rect 10798 1538 10958 8262
rect 12499 1538 12659 8262
rect 14200 1538 14360 8262
<< labels >>
rlabel metal2 s 14784 9600 14840 9900 6 bfg_out
port 1 nsew signal output
rlabel metal2 s 6048 100 6104 400 6 gf_out
port 2 nsew signal output
rlabel metal3 s 14600 3696 14900 3752 6 i0
port 3 nsew signal input
rlabel metal3 s 100 6048 400 6104 6 i1
port 4 nsew signal input
rlabel metal2 s 0 100 56 400 6 i2
port 5 nsew signal input
rlabel metal2 s 2352 9600 2408 9900 6 i3
port 6 nsew signal input
rlabel metal2 s 8736 9600 8792 9900 6 s0
port 7 nsew signal input
rlabel metal2 s 12432 100 12488 400 6 s1
port 8 nsew signal input
rlabel metal4 s 2293 1538 2453 8262 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 5695 1538 5855 8262 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 9097 1538 9257 8262 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 12499 1538 12659 8262 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 3994 1538 4154 8262 6 vss
port 10 nsew ground bidirectional
rlabel metal4 s 7396 1538 7556 8262 6 vss
port 10 nsew ground bidirectional
rlabel metal4 s 10798 1538 10958 8262 6 vss
port 10 nsew ground bidirectional
rlabel metal4 s 14200 1538 14360 8262 6 vss
port 10 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 187710
string GDS_FILE /home/aryap/src/bfg_mux_test_gf180mcu/openlane/bfg_mux_test_small/runs/22_12_12_00_59/results/signoff/bfg_mux_test_small.magic.gds
string GDS_START 77282
<< end >>

