(* blackbox *)
module gf180mcu_mux(
  input i0,
  input i1,
  input i2,
  input i3,
  input s0,
  input s0b,
  input s1,
  input s1b,
  output z
);
endmodule
