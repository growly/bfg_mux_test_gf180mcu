VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bfg_mux_test_small
  CLASS BLOCK ;
  FOREIGN bfg_mux_test_small ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 100.000 ;
  PIN bfg_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 96.000 148.400 99.000 ;
    END
  END bfg_out
  PIN gf_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 1.000 61.040 4.000 ;
    END
  END gf_out
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 146.000 36.960 149.000 37.520 ;
    END
  END i0
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 60.480 4.000 61.040 ;
    END
  END i1
  PIN i2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END i2
  PIN i3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 96.000 24.080 99.000 ;
    END
  END i3
  PIN s0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 96.000 87.920 99.000 ;
    END
  END s0
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1.000 124.880 4.000 ;
    END
  END s1
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.930 15.380 24.530 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 56.950 15.380 58.550 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 90.970 15.380 92.570 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 124.990 15.380 126.590 82.620 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 39.940 15.380 41.540 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 73.960 15.380 75.560 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 107.980 15.380 109.580 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 142.000 15.380 143.600 82.620 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 143.600 82.620 ;
      LAYER Metal2 ;
        RECT 0.140 95.700 23.220 96.000 ;
        RECT 24.380 95.700 87.060 96.000 ;
        RECT 88.220 95.700 147.540 96.000 ;
        RECT 0.140 4.300 148.260 95.700 ;
        RECT 0.860 4.000 60.180 4.300 ;
        RECT 61.340 4.000 124.020 4.300 ;
        RECT 125.180 4.000 148.260 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 61.340 148.310 88.900 ;
        RECT 0.090 60.180 0.700 61.340 ;
        RECT 4.300 60.180 148.310 61.340 ;
        RECT 0.090 37.820 148.310 60.180 ;
        RECT 0.090 36.660 145.700 37.820 ;
        RECT 0.090 12.460 148.310 36.660 ;
  END
END bfg_mux_test_small
END LIBRARY

