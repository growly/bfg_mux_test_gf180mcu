// This is the unpowered netlist.
module bfg_mux_test_small (bfg_out,
    gf_out,
    i0,
    i1,
    i2,
    i3,
    s0,
    s1);
 output bfg_out;
 output gf_out;
 input i0;
 input i1;
 input i2;
 input i3;
 input s0;
 input s1;

 wire _0_;
 wire _1_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2_ (.I(net5),
    .ZN(_0_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3_ (.I(net6),
    .ZN(_1_));
 gf180mcu_mux bfg_mux (.s0(net5),
    .z(net7),
    .i0_r(net1),
    .i2_r(net3),
    .i1_l(net2),
    .s0b(_0_),
    .i3_l(net4),
    .i0_l(net1),
    .i2_l(net3),
    .i1_r(net2),
    .s1b(_1_),
    .i3_r(net4),
    .s1(net6));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 gf_mux (.I0(net1),
    .I1(net2),
    .I2(net3),
    .I3(net4),
    .S0(net5),
    .S1(net6),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_80 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_81 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_82 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_83 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_84 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(i0),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(i1),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(i2),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(i3),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input5 (.I(s0),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(s1),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(bfg_out));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output8 (.I(net8),
    .Z(gf_out));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_s1b (.I(_1_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(i0));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(i1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(i2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(i3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(s0));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(s1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_gf_mux_I0 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_i0_l (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_i0_r (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_gf_mux_I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_i1_r (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_i1_l (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_gf_mux_I2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_i2_l (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_i2_r (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_gf_mux_I3 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_i3_r (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_i3_l (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_gf_mux_S0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_s0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_gf_mux_S1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_s1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bfg_mux_z (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_239 ();
endmodule

