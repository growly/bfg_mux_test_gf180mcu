magic
tech gf180mcuC
magscale 1 10
timestamp 1670835586
<< metal1 >>
rect 1344 16490 28560 16524
rect 1344 16438 4616 16490
rect 4668 16438 4720 16490
rect 4772 16438 4824 16490
rect 4876 16438 11420 16490
rect 11472 16438 11524 16490
rect 11576 16438 11628 16490
rect 11680 16438 18224 16490
rect 18276 16438 18328 16490
rect 18380 16438 18432 16490
rect 18484 16438 25028 16490
rect 25080 16438 25132 16490
rect 25184 16438 25236 16490
rect 25288 16438 28560 16490
rect 1344 16404 28560 16438
rect 4958 16210 5010 16222
rect 16830 16210 16882 16222
rect 7186 16158 7198 16210
rect 7250 16158 7262 16210
rect 26450 16158 26462 16210
rect 26514 16158 26526 16210
rect 4958 16146 5010 16158
rect 16830 16146 16882 16158
rect 25330 16046 25342 16098
rect 25394 16046 25406 16098
rect 5842 15934 5854 15986
rect 5906 15934 5918 15986
rect 19730 15934 19742 15986
rect 19794 15934 19806 15986
rect 17614 15874 17666 15886
rect 17614 15810 17666 15822
rect 24558 15874 24610 15886
rect 24558 15810 24610 15822
rect 1344 15706 28720 15740
rect 1344 15654 8018 15706
rect 8070 15654 8122 15706
rect 8174 15654 8226 15706
rect 8278 15654 14822 15706
rect 14874 15654 14926 15706
rect 14978 15654 15030 15706
rect 15082 15654 21626 15706
rect 21678 15654 21730 15706
rect 21782 15654 21834 15706
rect 21886 15654 28430 15706
rect 28482 15654 28534 15706
rect 28586 15654 28638 15706
rect 28690 15654 28720 15706
rect 1344 15620 28720 15654
rect 1344 14922 28560 14956
rect 1344 14870 4616 14922
rect 4668 14870 4720 14922
rect 4772 14870 4824 14922
rect 4876 14870 11420 14922
rect 11472 14870 11524 14922
rect 11576 14870 11628 14922
rect 11680 14870 18224 14922
rect 18276 14870 18328 14922
rect 18380 14870 18432 14922
rect 18484 14870 25028 14922
rect 25080 14870 25132 14922
rect 25184 14870 25236 14922
rect 25288 14870 28560 14922
rect 1344 14836 28560 14870
rect 1344 14138 28720 14172
rect 1344 14086 8018 14138
rect 8070 14086 8122 14138
rect 8174 14086 8226 14138
rect 8278 14086 14822 14138
rect 14874 14086 14926 14138
rect 14978 14086 15030 14138
rect 15082 14086 21626 14138
rect 21678 14086 21730 14138
rect 21782 14086 21834 14138
rect 21886 14086 28430 14138
rect 28482 14086 28534 14138
rect 28586 14086 28638 14138
rect 28690 14086 28720 14138
rect 1344 14052 28720 14086
rect 17614 13970 17666 13982
rect 17614 13906 17666 13918
rect 16606 13858 16658 13870
rect 16606 13794 16658 13806
rect 16494 13522 16546 13534
rect 16494 13458 16546 13470
rect 1344 13354 28560 13388
rect 1344 13302 4616 13354
rect 4668 13302 4720 13354
rect 4772 13302 4824 13354
rect 4876 13302 11420 13354
rect 11472 13302 11524 13354
rect 11576 13302 11628 13354
rect 11680 13302 18224 13354
rect 18276 13302 18328 13354
rect 18380 13302 18432 13354
rect 18484 13302 25028 13354
rect 25080 13302 25132 13354
rect 25184 13302 25236 13354
rect 25288 13302 28560 13354
rect 1344 13268 28560 13302
rect 3266 13022 3278 13074
rect 3330 13022 3342 13074
rect 7086 12850 7138 12862
rect 1922 12798 1934 12850
rect 1986 12798 1998 12850
rect 7086 12786 7138 12798
rect 7646 12850 7698 12862
rect 7646 12786 7698 12798
rect 7198 12738 7250 12750
rect 7198 12674 7250 12686
rect 1344 12570 28720 12604
rect 1344 12518 8018 12570
rect 8070 12518 8122 12570
rect 8174 12518 8226 12570
rect 8278 12518 14822 12570
rect 14874 12518 14926 12570
rect 14978 12518 15030 12570
rect 15082 12518 21626 12570
rect 21678 12518 21730 12570
rect 21782 12518 21834 12570
rect 21886 12518 28430 12570
rect 28482 12518 28534 12570
rect 28586 12518 28638 12570
rect 28690 12518 28720 12570
rect 1344 12484 28720 12518
rect 1710 12178 1762 12190
rect 1710 12114 1762 12126
rect 1344 11786 28560 11820
rect 1344 11734 4616 11786
rect 4668 11734 4720 11786
rect 4772 11734 4824 11786
rect 4876 11734 11420 11786
rect 11472 11734 11524 11786
rect 11576 11734 11628 11786
rect 11680 11734 18224 11786
rect 18276 11734 18328 11786
rect 18380 11734 18432 11786
rect 18484 11734 25028 11786
rect 25080 11734 25132 11786
rect 25184 11734 25236 11786
rect 25288 11734 28560 11786
rect 1344 11700 28560 11734
rect 12798 11506 12850 11518
rect 12798 11442 12850 11454
rect 13582 11506 13634 11518
rect 13582 11442 13634 11454
rect 14142 11506 14194 11518
rect 14142 11442 14194 11454
rect 14478 11506 14530 11518
rect 14478 11442 14530 11454
rect 15262 11506 15314 11518
rect 15262 11442 15314 11454
rect 15710 11506 15762 11518
rect 15710 11442 15762 11454
rect 1344 11002 28720 11036
rect 1344 10950 8018 11002
rect 8070 10950 8122 11002
rect 8174 10950 8226 11002
rect 8278 10950 14822 11002
rect 14874 10950 14926 11002
rect 14978 10950 15030 11002
rect 15082 10950 21626 11002
rect 21678 10950 21730 11002
rect 21782 10950 21834 11002
rect 21886 10950 28430 11002
rect 28482 10950 28534 11002
rect 28586 10950 28638 11002
rect 28690 10950 28720 11002
rect 1344 10916 28720 10950
rect 15138 10782 15150 10834
rect 15202 10831 15214 10834
rect 15698 10831 15710 10834
rect 15202 10785 15710 10831
rect 15202 10782 15214 10785
rect 15698 10782 15710 10785
rect 15762 10782 15774 10834
rect 1344 10218 10976 10252
rect 1344 10166 4616 10218
rect 4668 10166 4720 10218
rect 4772 10166 4824 10218
rect 4876 10166 10976 10218
rect 1344 10132 10976 10166
rect 17808 10218 28560 10252
rect 17808 10166 18224 10218
rect 18276 10166 18328 10218
rect 18380 10166 18432 10218
rect 18484 10166 25028 10218
rect 25080 10166 25132 10218
rect 25184 10166 25236 10218
rect 25288 10166 28560 10218
rect 17808 10132 28560 10166
rect 1344 9434 10976 9468
rect 1344 9382 8018 9434
rect 8070 9382 8122 9434
rect 8174 9382 8226 9434
rect 8278 9382 10976 9434
rect 1344 9348 10976 9382
rect 17808 9434 28720 9468
rect 17808 9382 21626 9434
rect 21678 9382 21730 9434
rect 21782 9382 21834 9434
rect 21886 9382 28430 9434
rect 28482 9382 28534 9434
rect 28586 9382 28638 9434
rect 28690 9382 28720 9434
rect 15250 9375 15262 9378
rect 13473 9329 15262 9375
rect 10110 8930 10162 8942
rect 10110 8866 10162 8878
rect 10558 8930 10610 8942
rect 10558 8866 10610 8878
rect 1344 8650 10976 8684
rect 1344 8598 4616 8650
rect 4668 8598 4720 8650
rect 4772 8598 4824 8650
rect 4876 8598 10976 8650
rect 13473 8608 13519 9329
rect 15250 9326 15262 9329
rect 15314 9326 15326 9378
rect 17808 9348 28720 9382
rect 13570 9214 13582 9266
rect 13634 9263 13646 9266
rect 13634 9217 14243 9263
rect 13634 9214 13646 9217
rect 14018 9039 14030 9042
rect 13865 8993 14030 9039
rect 13865 8613 13911 8993
rect 14018 8990 14030 8993
rect 14082 8990 14094 9042
rect 14197 8733 14243 9217
rect 18286 8930 18338 8942
rect 18286 8866 18338 8878
rect 18622 8930 18674 8942
rect 18622 8866 18674 8878
rect 15026 8815 15038 8818
rect 14929 8769 15038 8815
rect 1344 8564 10976 8598
rect 14130 8573 14142 8625
rect 14194 8573 14206 8625
rect 14929 8581 14975 8769
rect 15026 8766 15038 8769
rect 15090 8766 15102 8818
rect 15250 8606 15262 8658
rect 15314 8606 15326 8658
rect 17808 8650 28560 8684
rect 17808 8598 18224 8650
rect 18276 8598 18328 8650
rect 18380 8598 18432 8650
rect 18484 8598 25028 8650
rect 25080 8598 25132 8650
rect 25184 8598 25236 8650
rect 25288 8598 28560 8650
rect 17808 8564 28560 8598
rect 13090 8407 13102 8459
rect 13154 8407 13166 8459
rect 15452 8430 15464 8482
rect 15516 8430 15528 8482
rect 24882 8318 24894 8370
rect 24946 8318 24958 8370
rect 13090 8244 13102 8296
rect 13154 8244 13166 8296
rect 15457 8248 15469 8300
rect 15521 8248 15533 8300
rect 18174 8146 18226 8158
rect 12786 8069 12798 8121
rect 12850 8118 12862 8121
rect 12850 8072 13160 8118
rect 12850 8069 12862 8072
rect 14914 8069 14926 8121
rect 14978 8118 14990 8121
rect 14978 8072 15064 8118
rect 26226 8094 26238 8146
rect 26290 8094 26302 8146
rect 18174 8082 18226 8094
rect 14978 8069 14990 8072
rect 10446 8034 10498 8046
rect 14435 8031 14481 8051
rect 26910 8034 26962 8046
rect 14578 8031 14590 8034
rect 14435 7985 14590 8031
rect 14578 7982 14590 7985
rect 14642 7982 14654 8034
rect 10446 7970 10498 7982
rect 26910 7970 26962 7982
rect 1344 7866 10976 7900
rect 1344 7814 8018 7866
rect 8070 7814 8122 7866
rect 8174 7814 8226 7866
rect 8278 7814 10976 7866
rect 1344 7780 10976 7814
rect 17808 7866 28720 7900
rect 17808 7814 21626 7866
rect 21678 7814 21730 7866
rect 21782 7814 21834 7866
rect 21886 7814 28430 7866
rect 28482 7814 28534 7866
rect 28586 7814 28638 7866
rect 28690 7814 28720 7866
rect 17808 7780 28720 7814
rect 1344 7082 10976 7116
rect 1344 7030 4616 7082
rect 4668 7030 4720 7082
rect 4772 7030 4824 7082
rect 4876 7030 10976 7082
rect 1344 6996 10976 7030
rect 17808 7082 28560 7116
rect 17808 7030 18224 7082
rect 18276 7030 18328 7082
rect 18380 7030 18432 7082
rect 18484 7030 25028 7082
rect 25080 7030 25132 7082
rect 25184 7030 25236 7082
rect 25288 7030 28560 7082
rect 17808 6996 28560 7030
rect 1344 6298 10976 6332
rect 1344 6246 8018 6298
rect 8070 6246 8122 6298
rect 8174 6246 8226 6298
rect 8278 6246 10976 6298
rect 1344 6212 10976 6246
rect 17808 6298 28720 6332
rect 17808 6246 21626 6298
rect 21678 6246 21730 6298
rect 21782 6246 21834 6298
rect 21886 6246 28430 6298
rect 28482 6246 28534 6298
rect 28586 6246 28638 6298
rect 28690 6246 28720 6298
rect 17808 6212 28720 6246
rect 1344 5514 28560 5548
rect 1344 5462 4616 5514
rect 4668 5462 4720 5514
rect 4772 5462 4824 5514
rect 4876 5462 11420 5514
rect 11472 5462 11524 5514
rect 11576 5462 11628 5514
rect 11680 5462 18224 5514
rect 18276 5462 18328 5514
rect 18380 5462 18432 5514
rect 18484 5462 25028 5514
rect 25080 5462 25132 5514
rect 25184 5462 25236 5514
rect 25288 5462 28560 5514
rect 1344 5428 28560 5462
rect 1344 4730 28720 4764
rect 1344 4678 8018 4730
rect 8070 4678 8122 4730
rect 8174 4678 8226 4730
rect 8278 4678 14822 4730
rect 14874 4678 14926 4730
rect 14978 4678 15030 4730
rect 15082 4678 21626 4730
rect 21678 4678 21730 4730
rect 21782 4678 21834 4730
rect 21886 4678 28430 4730
rect 28482 4678 28534 4730
rect 28586 4678 28638 4730
rect 28690 4678 28720 4730
rect 1344 4644 28720 4678
rect 3278 4562 3330 4574
rect 3278 4498 3330 4510
rect 3614 4562 3666 4574
rect 3614 4498 3666 4510
rect 7870 4562 7922 4574
rect 7870 4498 7922 4510
rect 8766 4562 8818 4574
rect 8766 4498 8818 4510
rect 7422 4450 7474 4462
rect 6402 4398 6414 4450
rect 6466 4398 6478 4450
rect 7422 4386 7474 4398
rect 5966 4338 6018 4350
rect 8318 4338 8370 4350
rect 4386 4286 4398 4338
rect 4450 4286 4462 4338
rect 5170 4286 5182 4338
rect 5234 4286 5246 4338
rect 6626 4286 6638 4338
rect 6690 4286 6702 4338
rect 7074 4286 7086 4338
rect 7138 4286 7150 4338
rect 5966 4274 6018 4286
rect 8318 4274 8370 4286
rect 1822 4226 1874 4238
rect 1822 4162 1874 4174
rect 1344 3946 28560 3980
rect 1344 3894 4616 3946
rect 4668 3894 4720 3946
rect 4772 3894 4824 3946
rect 4876 3894 11420 3946
rect 11472 3894 11524 3946
rect 11576 3894 11628 3946
rect 11680 3894 18224 3946
rect 18276 3894 18328 3946
rect 18380 3894 18432 3946
rect 18484 3894 25028 3946
rect 25080 3894 25132 3946
rect 25184 3894 25236 3946
rect 25288 3894 28560 3946
rect 1344 3860 28560 3894
rect 7758 3666 7810 3678
rect 3266 3614 3278 3666
rect 3330 3614 3342 3666
rect 12226 3614 12238 3666
rect 12290 3614 12302 3666
rect 25330 3614 25342 3666
rect 25394 3614 25406 3666
rect 7758 3602 7810 3614
rect 11554 3502 11566 3554
rect 11618 3502 11630 3554
rect 24670 3442 24722 3454
rect 1922 3390 1934 3442
rect 1986 3390 1998 3442
rect 26338 3390 26350 3442
rect 26402 3390 26414 3442
rect 24670 3378 24722 3390
rect 1344 3162 28720 3196
rect 1344 3110 8018 3162
rect 8070 3110 8122 3162
rect 8174 3110 8226 3162
rect 8278 3110 14822 3162
rect 14874 3110 14926 3162
rect 14978 3110 15030 3162
rect 15082 3110 21626 3162
rect 21678 3110 21730 3162
rect 21782 3110 21834 3162
rect 21886 3110 28430 3162
rect 28482 3110 28534 3162
rect 28586 3110 28638 3162
rect 28690 3110 28720 3162
rect 1344 3076 28720 3110
<< via1 >>
rect 4616 16438 4668 16490
rect 4720 16438 4772 16490
rect 4824 16438 4876 16490
rect 11420 16438 11472 16490
rect 11524 16438 11576 16490
rect 11628 16438 11680 16490
rect 18224 16438 18276 16490
rect 18328 16438 18380 16490
rect 18432 16438 18484 16490
rect 25028 16438 25080 16490
rect 25132 16438 25184 16490
rect 25236 16438 25288 16490
rect 4958 16158 5010 16210
rect 7198 16158 7250 16210
rect 16830 16158 16882 16210
rect 26462 16158 26514 16210
rect 25342 16046 25394 16098
rect 5854 15934 5906 15986
rect 19742 15934 19794 15986
rect 17614 15822 17666 15874
rect 24558 15822 24610 15874
rect 8018 15654 8070 15706
rect 8122 15654 8174 15706
rect 8226 15654 8278 15706
rect 14822 15654 14874 15706
rect 14926 15654 14978 15706
rect 15030 15654 15082 15706
rect 21626 15654 21678 15706
rect 21730 15654 21782 15706
rect 21834 15654 21886 15706
rect 28430 15654 28482 15706
rect 28534 15654 28586 15706
rect 28638 15654 28690 15706
rect 4616 14870 4668 14922
rect 4720 14870 4772 14922
rect 4824 14870 4876 14922
rect 11420 14870 11472 14922
rect 11524 14870 11576 14922
rect 11628 14870 11680 14922
rect 18224 14870 18276 14922
rect 18328 14870 18380 14922
rect 18432 14870 18484 14922
rect 25028 14870 25080 14922
rect 25132 14870 25184 14922
rect 25236 14870 25288 14922
rect 8018 14086 8070 14138
rect 8122 14086 8174 14138
rect 8226 14086 8278 14138
rect 14822 14086 14874 14138
rect 14926 14086 14978 14138
rect 15030 14086 15082 14138
rect 21626 14086 21678 14138
rect 21730 14086 21782 14138
rect 21834 14086 21886 14138
rect 28430 14086 28482 14138
rect 28534 14086 28586 14138
rect 28638 14086 28690 14138
rect 17614 13918 17666 13970
rect 16606 13806 16658 13858
rect 16494 13470 16546 13522
rect 4616 13302 4668 13354
rect 4720 13302 4772 13354
rect 4824 13302 4876 13354
rect 11420 13302 11472 13354
rect 11524 13302 11576 13354
rect 11628 13302 11680 13354
rect 18224 13302 18276 13354
rect 18328 13302 18380 13354
rect 18432 13302 18484 13354
rect 25028 13302 25080 13354
rect 25132 13302 25184 13354
rect 25236 13302 25288 13354
rect 3278 13022 3330 13074
rect 1934 12798 1986 12850
rect 7086 12798 7138 12850
rect 7646 12798 7698 12850
rect 7198 12686 7250 12738
rect 8018 12518 8070 12570
rect 8122 12518 8174 12570
rect 8226 12518 8278 12570
rect 14822 12518 14874 12570
rect 14926 12518 14978 12570
rect 15030 12518 15082 12570
rect 21626 12518 21678 12570
rect 21730 12518 21782 12570
rect 21834 12518 21886 12570
rect 28430 12518 28482 12570
rect 28534 12518 28586 12570
rect 28638 12518 28690 12570
rect 1710 12126 1762 12178
rect 4616 11734 4668 11786
rect 4720 11734 4772 11786
rect 4824 11734 4876 11786
rect 11420 11734 11472 11786
rect 11524 11734 11576 11786
rect 11628 11734 11680 11786
rect 18224 11734 18276 11786
rect 18328 11734 18380 11786
rect 18432 11734 18484 11786
rect 25028 11734 25080 11786
rect 25132 11734 25184 11786
rect 25236 11734 25288 11786
rect 12798 11454 12850 11506
rect 13582 11454 13634 11506
rect 14142 11454 14194 11506
rect 14478 11454 14530 11506
rect 15262 11454 15314 11506
rect 15710 11454 15762 11506
rect 8018 10950 8070 11002
rect 8122 10950 8174 11002
rect 8226 10950 8278 11002
rect 14822 10950 14874 11002
rect 14926 10950 14978 11002
rect 15030 10950 15082 11002
rect 21626 10950 21678 11002
rect 21730 10950 21782 11002
rect 21834 10950 21886 11002
rect 28430 10950 28482 11002
rect 28534 10950 28586 11002
rect 28638 10950 28690 11002
rect 15150 10782 15202 10834
rect 15710 10782 15762 10834
rect 4616 10166 4668 10218
rect 4720 10166 4772 10218
rect 4824 10166 4876 10218
rect 18224 10166 18276 10218
rect 18328 10166 18380 10218
rect 18432 10166 18484 10218
rect 25028 10166 25080 10218
rect 25132 10166 25184 10218
rect 25236 10166 25288 10218
rect 8018 9382 8070 9434
rect 8122 9382 8174 9434
rect 8226 9382 8278 9434
rect 21626 9382 21678 9434
rect 21730 9382 21782 9434
rect 21834 9382 21886 9434
rect 28430 9382 28482 9434
rect 28534 9382 28586 9434
rect 28638 9382 28690 9434
rect 10110 8878 10162 8930
rect 10558 8878 10610 8930
rect 4616 8598 4668 8650
rect 4720 8598 4772 8650
rect 4824 8598 4876 8650
rect 15262 9326 15314 9378
rect 13582 9214 13634 9266
rect 14030 8990 14082 9042
rect 18286 8878 18338 8930
rect 18622 8878 18674 8930
rect 14142 8573 14194 8625
rect 15038 8766 15090 8818
rect 15262 8606 15314 8658
rect 18224 8598 18276 8650
rect 18328 8598 18380 8650
rect 18432 8598 18484 8650
rect 25028 8598 25080 8650
rect 25132 8598 25184 8650
rect 25236 8598 25288 8650
rect 13102 8407 13154 8459
rect 15464 8430 15516 8482
rect 24894 8318 24946 8370
rect 13102 8244 13154 8296
rect 15469 8248 15521 8300
rect 12798 8069 12850 8121
rect 14926 8069 14978 8121
rect 18174 8094 18226 8146
rect 26238 8094 26290 8146
rect 10446 7982 10498 8034
rect 14590 7982 14642 8034
rect 26910 7982 26962 8034
rect 8018 7814 8070 7866
rect 8122 7814 8174 7866
rect 8226 7814 8278 7866
rect 21626 7814 21678 7866
rect 21730 7814 21782 7866
rect 21834 7814 21886 7866
rect 28430 7814 28482 7866
rect 28534 7814 28586 7866
rect 28638 7814 28690 7866
rect 4616 7030 4668 7082
rect 4720 7030 4772 7082
rect 4824 7030 4876 7082
rect 18224 7030 18276 7082
rect 18328 7030 18380 7082
rect 18432 7030 18484 7082
rect 25028 7030 25080 7082
rect 25132 7030 25184 7082
rect 25236 7030 25288 7082
rect 8018 6246 8070 6298
rect 8122 6246 8174 6298
rect 8226 6246 8278 6298
rect 21626 6246 21678 6298
rect 21730 6246 21782 6298
rect 21834 6246 21886 6298
rect 28430 6246 28482 6298
rect 28534 6246 28586 6298
rect 28638 6246 28690 6298
rect 4616 5462 4668 5514
rect 4720 5462 4772 5514
rect 4824 5462 4876 5514
rect 11420 5462 11472 5514
rect 11524 5462 11576 5514
rect 11628 5462 11680 5514
rect 18224 5462 18276 5514
rect 18328 5462 18380 5514
rect 18432 5462 18484 5514
rect 25028 5462 25080 5514
rect 25132 5462 25184 5514
rect 25236 5462 25288 5514
rect 8018 4678 8070 4730
rect 8122 4678 8174 4730
rect 8226 4678 8278 4730
rect 14822 4678 14874 4730
rect 14926 4678 14978 4730
rect 15030 4678 15082 4730
rect 21626 4678 21678 4730
rect 21730 4678 21782 4730
rect 21834 4678 21886 4730
rect 28430 4678 28482 4730
rect 28534 4678 28586 4730
rect 28638 4678 28690 4730
rect 3278 4510 3330 4562
rect 3614 4510 3666 4562
rect 7870 4510 7922 4562
rect 8766 4510 8818 4562
rect 6414 4398 6466 4450
rect 7422 4398 7474 4450
rect 4398 4286 4450 4338
rect 5182 4286 5234 4338
rect 5966 4286 6018 4338
rect 6638 4286 6690 4338
rect 7086 4286 7138 4338
rect 8318 4286 8370 4338
rect 1822 4174 1874 4226
rect 4616 3894 4668 3946
rect 4720 3894 4772 3946
rect 4824 3894 4876 3946
rect 11420 3894 11472 3946
rect 11524 3894 11576 3946
rect 11628 3894 11680 3946
rect 18224 3894 18276 3946
rect 18328 3894 18380 3946
rect 18432 3894 18484 3946
rect 25028 3894 25080 3946
rect 25132 3894 25184 3946
rect 25236 3894 25288 3946
rect 3278 3614 3330 3666
rect 7758 3614 7810 3666
rect 12238 3614 12290 3666
rect 25342 3614 25394 3666
rect 11566 3502 11618 3554
rect 1934 3390 1986 3442
rect 24670 3390 24722 3442
rect 26350 3390 26402 3442
rect 8018 3110 8070 3162
rect 8122 3110 8174 3162
rect 8226 3110 8278 3162
rect 14822 3110 14874 3162
rect 14926 3110 14978 3162
rect 15030 3110 15082 3162
rect 21626 3110 21678 3162
rect 21730 3110 21782 3162
rect 21834 3110 21886 3162
rect 28430 3110 28482 3162
rect 28534 3110 28586 3162
rect 28638 3110 28690 3162
<< metal2 >>
rect 4704 19200 4816 19800
rect 17472 19200 17584 19800
rect 29568 19200 29680 19800
rect 4732 17108 4788 19200
rect 4732 17052 5012 17108
rect 4614 16492 4878 16502
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4614 16426 4878 16436
rect 4956 16210 5012 17052
rect 11418 16492 11682 16502
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11418 16426 11682 16436
rect 4956 16158 4958 16210
rect 5010 16158 5012 16210
rect 4956 15988 5012 16158
rect 7196 16212 7252 16222
rect 7196 16118 7252 16156
rect 10444 16212 10500 16222
rect 4956 15922 5012 15932
rect 5852 15988 5908 15998
rect 5852 15894 5908 15932
rect 8016 15708 8280 15718
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8016 15642 8280 15652
rect 4614 14924 4878 14934
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4614 14858 4878 14868
rect 8016 14140 8280 14150
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8016 14074 8280 14084
rect 4614 13356 4878 13366
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4614 13290 4878 13300
rect 3276 13076 3332 13086
rect 3276 13074 3444 13076
rect 3276 13022 3278 13074
rect 3330 13022 3444 13074
rect 3276 13020 3444 13022
rect 3276 13010 3332 13020
rect 1932 12852 1988 12862
rect 1708 12850 1988 12852
rect 1708 12798 1934 12850
rect 1986 12798 1988 12850
rect 1708 12796 1988 12798
rect 1708 12180 1764 12796
rect 1932 12786 1988 12796
rect 1708 12086 1764 12124
rect 3388 11956 3444 13020
rect 7084 12852 7140 12862
rect 7084 12758 7140 12796
rect 7644 12852 7700 12862
rect 7644 12758 7700 12796
rect 7196 12740 7252 12750
rect 7196 12646 7252 12684
rect 8016 12572 8280 12582
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8016 12506 8280 12516
rect 3388 11890 3444 11900
rect 3612 11956 3668 11966
rect 3276 4564 3332 4574
rect 1820 4228 1876 4238
rect 1820 4226 1988 4228
rect 1820 4174 1822 4226
rect 1874 4174 1988 4226
rect 1820 4172 1988 4174
rect 1820 4162 1876 4172
rect 1932 3442 1988 4172
rect 3276 3666 3332 4508
rect 3612 4562 3668 11900
rect 4614 11788 4878 11798
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4614 11722 4878 11732
rect 8016 11004 8280 11014
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8016 10938 8280 10948
rect 4614 10220 4878 10230
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4614 10154 4878 10164
rect 8016 9436 8280 9446
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8016 9370 8280 9380
rect 7756 8932 7812 8942
rect 4614 8652 4878 8662
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4614 8586 4878 8596
rect 4614 7084 4878 7094
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4614 7018 4878 7028
rect 7420 6916 7476 6926
rect 4614 5516 4878 5526
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4614 5450 4878 5460
rect 3612 4510 3614 4562
rect 3666 4510 3668 4562
rect 3612 4340 3668 4510
rect 6748 4900 6804 4910
rect 3612 4274 3668 4284
rect 4396 4452 4452 4462
rect 4396 4338 4452 4396
rect 6412 4450 6468 4462
rect 6412 4398 6414 4450
rect 6466 4398 6468 4450
rect 4396 4286 4398 4338
rect 4450 4286 4452 4338
rect 4396 4274 4452 4286
rect 5180 4340 5236 4350
rect 5180 4246 5236 4284
rect 5964 4340 6020 4350
rect 5964 4246 6020 4284
rect 4614 3948 4878 3958
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4614 3882 4878 3892
rect 3276 3614 3278 3666
rect 3330 3614 3332 3666
rect 3276 3602 3332 3614
rect 6412 3556 6468 4398
rect 6636 4340 6692 4350
rect 6748 4340 6804 4844
rect 7420 4564 7476 6860
rect 7420 4450 7476 4508
rect 7420 4398 7422 4450
rect 7474 4398 7476 4450
rect 7420 4386 7476 4398
rect 7756 4452 7812 8876
rect 10108 8930 10164 8942
rect 10108 8878 10110 8930
rect 10162 8878 10164 8930
rect 10108 8260 10164 8878
rect 8016 7868 8280 7878
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8016 7802 8280 7812
rect 10108 6916 10164 8204
rect 10108 6850 10164 6860
rect 10444 8148 10500 16156
rect 16828 16212 16884 16222
rect 16828 16118 16884 16156
rect 17500 16212 17556 19200
rect 26460 17780 26516 17790
rect 18222 16492 18486 16502
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18222 16426 18486 16436
rect 25026 16492 25290 16502
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25026 16426 25290 16436
rect 17500 16146 17556 16156
rect 19740 16212 19796 16222
rect 19740 15986 19796 16156
rect 26460 16210 26516 17724
rect 29596 17780 29652 19200
rect 29596 17714 29652 17724
rect 26460 16158 26462 16210
rect 26514 16158 26516 16210
rect 26460 16146 26516 16158
rect 19740 15934 19742 15986
rect 19794 15934 19796 15986
rect 19740 15922 19796 15934
rect 25340 16098 25396 16110
rect 25340 16046 25342 16098
rect 25394 16046 25396 16098
rect 17612 15874 17668 15886
rect 17612 15822 17614 15874
rect 17666 15822 17668 15874
rect 14820 15708 15084 15718
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 14820 15642 15084 15652
rect 14140 15540 14196 15550
rect 11418 14924 11682 14934
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11418 14858 11682 14868
rect 14028 13524 14084 13534
rect 11418 13356 11682 13366
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11418 13290 11682 13300
rect 13580 12740 13636 12750
rect 12796 11956 12852 11966
rect 11418 11788 11682 11798
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11418 11722 11682 11732
rect 12796 11506 12852 11900
rect 12796 11454 12798 11506
rect 12850 11454 12852 11506
rect 12796 11442 12852 11454
rect 13580 11506 13636 12684
rect 13580 11454 13582 11506
rect 13634 11454 13636 11506
rect 13580 9266 13636 11454
rect 13580 9214 13582 9266
rect 13634 9214 13636 9266
rect 13580 9202 13636 9214
rect 14028 9042 14084 13468
rect 14028 8990 14030 9042
rect 14082 8990 14084 9042
rect 14028 8978 14084 8990
rect 14140 11506 14196 15484
rect 14820 14140 15084 14150
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 14820 14074 15084 14084
rect 17612 13970 17668 15822
rect 24556 15874 24612 15886
rect 24556 15822 24558 15874
rect 24610 15822 24612 15874
rect 21624 15708 21888 15718
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21624 15642 21888 15652
rect 24556 15540 24612 15822
rect 24556 15474 24612 15484
rect 25340 15540 25396 16046
rect 28428 15708 28692 15718
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28428 15642 28692 15652
rect 25340 15474 25396 15484
rect 18222 14924 18486 14934
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18222 14858 18486 14868
rect 25026 14924 25290 14934
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25026 14858 25290 14868
rect 21624 14140 21888 14150
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21624 14074 21888 14084
rect 28428 14140 28692 14150
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28428 14074 28692 14084
rect 17612 13918 17614 13970
rect 17666 13918 17668 13970
rect 15708 13860 15764 13870
rect 14140 11454 14142 11506
rect 14194 11454 14196 11506
rect 10556 8932 10612 8942
rect 10556 8484 10612 8876
rect 14140 8625 14196 11454
rect 14140 8573 14142 8625
rect 14194 8573 14196 8625
rect 14140 8561 14196 8573
rect 14476 12852 14532 12862
rect 14476 11506 14532 12796
rect 14820 12572 15084 12582
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 14820 12506 15084 12516
rect 14476 11454 14478 11506
rect 14530 11454 14532 11506
rect 10556 8418 10612 8428
rect 13100 8484 13156 8499
rect 13100 8407 13102 8428
rect 13154 8407 13156 8428
rect 13100 8395 13156 8407
rect 13100 8296 13156 8308
rect 13100 8260 13102 8296
rect 13154 8260 13156 8296
rect 13100 8194 13156 8204
rect 10444 8034 10500 8092
rect 12796 8148 12852 8158
rect 12796 8069 12798 8092
rect 12850 8069 12852 8092
rect 12796 8054 12852 8069
rect 10444 7982 10446 8034
rect 10498 7982 10500 8034
rect 8016 6300 8280 6310
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8016 6234 8280 6244
rect 7868 4900 7924 4910
rect 7868 4562 7924 4844
rect 10444 4900 10500 7982
rect 14476 8036 14532 11454
rect 15260 11956 15316 11966
rect 15260 11506 15316 11900
rect 15260 11454 15262 11506
rect 15314 11454 15316 11506
rect 14820 11004 15084 11014
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 14820 10938 15084 10948
rect 15148 10834 15204 10846
rect 15148 10782 15150 10834
rect 15202 10782 15204 10834
rect 15036 8820 15092 8830
rect 15148 8820 15204 10782
rect 15036 8818 15204 8820
rect 15036 8766 15038 8818
rect 15090 8766 15204 8818
rect 15036 8764 15204 8766
rect 15036 8754 15092 8764
rect 14924 8148 14980 8158
rect 14924 8069 14926 8092
rect 14978 8069 14980 8092
rect 14924 8054 14980 8069
rect 14588 8036 14644 8046
rect 14476 8034 14644 8036
rect 14476 7982 14590 8034
rect 14642 7982 14644 8034
rect 14476 7980 14644 7982
rect 11418 5516 11682 5526
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11418 5450 11682 5460
rect 10444 4834 10500 4844
rect 8016 4732 8280 4742
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8016 4666 8280 4676
rect 7868 4510 7870 4562
rect 7922 4510 7924 4562
rect 7868 4498 7924 4510
rect 8764 4564 8820 4574
rect 6636 4338 6804 4340
rect 6636 4286 6638 4338
rect 6690 4286 6804 4338
rect 6636 4284 6804 4286
rect 7084 4338 7140 4350
rect 7084 4286 7086 4338
rect 7138 4286 7140 4338
rect 6636 4274 6692 4284
rect 7084 4228 7140 4286
rect 7084 4162 7140 4172
rect 7756 3666 7812 4396
rect 8316 4340 8372 4350
rect 8316 4246 8372 4284
rect 8764 4228 8820 4508
rect 8764 4162 8820 4172
rect 14476 4340 14532 7980
rect 14588 7970 14644 7980
rect 14820 4732 15084 4742
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 14820 4666 15084 4676
rect 15148 4564 15204 8764
rect 15260 9378 15316 11454
rect 15708 11506 15764 13804
rect 16604 13860 16660 13870
rect 16604 13766 16660 13804
rect 17612 13860 17668 13918
rect 17612 13794 17668 13804
rect 16492 13524 16548 13534
rect 16492 13430 16548 13468
rect 18222 13356 18486 13366
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18222 13290 18486 13300
rect 25026 13356 25290 13366
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25026 13290 25290 13300
rect 21624 12572 21888 12582
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21624 12506 21888 12516
rect 28428 12572 28692 12582
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28428 12506 28692 12516
rect 18222 11788 18486 11798
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18222 11722 18486 11732
rect 25026 11788 25290 11798
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25026 11722 25290 11732
rect 15708 11454 15710 11506
rect 15762 11454 15764 11506
rect 15708 10834 15764 11454
rect 21624 11004 21888 11014
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21624 10938 21888 10948
rect 28428 11004 28692 11014
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28428 10938 28692 10948
rect 15708 10782 15710 10834
rect 15762 10782 15764 10834
rect 15708 10770 15764 10782
rect 18222 10220 18486 10230
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18222 10154 18486 10164
rect 25026 10220 25290 10230
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25026 10154 25290 10164
rect 15260 9326 15262 9378
rect 15314 9326 15316 9378
rect 21624 9436 21888 9446
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21624 9370 21888 9380
rect 28428 9436 28692 9446
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28428 9370 28692 9380
rect 15260 8658 15316 9326
rect 18284 8932 18340 8942
rect 15260 8606 15262 8658
rect 15314 8606 15316 8658
rect 15260 8594 15316 8606
rect 18060 8930 18340 8932
rect 18060 8878 18286 8930
rect 18338 8878 18340 8930
rect 18060 8876 18340 8878
rect 15462 8484 15518 8522
rect 15462 8418 15518 8428
rect 18060 8484 18116 8876
rect 18284 8820 18340 8876
rect 18284 8754 18340 8764
rect 18620 8930 18676 8942
rect 18620 8878 18622 8930
rect 18674 8878 18676 8930
rect 18222 8652 18486 8662
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18222 8586 18486 8596
rect 18060 8418 18116 8428
rect 15467 8300 15523 8312
rect 15467 8260 15469 8300
rect 15521 8260 15523 8300
rect 15467 8194 15523 8204
rect 18620 8260 18676 8878
rect 24892 8820 24948 8830
rect 24892 8370 24948 8764
rect 25026 8652 25290 8662
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25026 8586 25290 8596
rect 24892 8318 24894 8370
rect 24946 8318 24948 8370
rect 24892 8306 24948 8318
rect 18620 8194 18676 8204
rect 18172 8148 18228 8158
rect 18172 8054 18228 8092
rect 26236 8148 26292 8158
rect 26236 8054 26292 8092
rect 26908 8148 26964 8158
rect 26908 8034 26964 8092
rect 26908 7982 26910 8034
rect 26962 7982 26964 8034
rect 21624 7868 21888 7878
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21624 7802 21888 7812
rect 26908 7476 26964 7982
rect 28428 7868 28692 7878
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28428 7802 28692 7812
rect 26908 7410 26964 7420
rect 18222 7084 18486 7094
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18222 7018 18486 7028
rect 25026 7084 25290 7094
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25026 7018 25290 7028
rect 21624 6300 21888 6310
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21624 6234 21888 6244
rect 28428 6300 28692 6310
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28428 6234 28692 6244
rect 18222 5516 18486 5526
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18222 5450 18486 5460
rect 25026 5516 25290 5526
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25026 5450 25290 5460
rect 21624 4732 21888 4742
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21624 4666 21888 4676
rect 28428 4732 28692 4742
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28428 4666 28692 4676
rect 15148 4498 15204 4508
rect 11418 3948 11682 3958
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11418 3882 11682 3892
rect 12236 3668 12292 3678
rect 7756 3614 7758 3666
rect 7810 3614 7812 3666
rect 7756 3602 7812 3614
rect 12124 3666 12292 3668
rect 12124 3614 12238 3666
rect 12290 3614 12292 3666
rect 12124 3612 12292 3614
rect 6412 3490 6468 3500
rect 11564 3556 11620 3566
rect 11564 3462 11620 3500
rect 1932 3390 1934 3442
rect 1986 3390 1988 3442
rect 28 2548 84 2558
rect 28 800 84 2492
rect 1932 2548 1988 3390
rect 8016 3164 8280 3174
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8016 3098 8280 3108
rect 1932 2482 1988 2492
rect 12124 800 12180 3612
rect 12236 3602 12292 3612
rect 14476 3668 14532 4284
rect 18222 3948 18486 3958
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18222 3882 18486 3892
rect 25026 3948 25290 3958
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25026 3882 25290 3892
rect 14476 3602 14532 3612
rect 25340 3668 25396 3678
rect 25340 3574 25396 3612
rect 24668 3444 24724 3454
rect 24892 3444 24948 3454
rect 24668 3442 24892 3444
rect 24668 3390 24670 3442
rect 24722 3390 24892 3442
rect 24668 3388 24892 3390
rect 24668 3378 24724 3388
rect 14820 3164 15084 3174
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 14820 3098 15084 3108
rect 21624 3164 21888 3174
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21624 3098 21888 3108
rect 24892 800 24948 3388
rect 26348 3444 26404 3454
rect 26348 3350 26404 3388
rect 28428 3164 28692 3174
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28428 3098 28692 3108
rect 0 200 112 800
rect 12096 200 12208 800
rect 24864 200 24976 800
<< via2 >>
rect 4614 16490 4670 16492
rect 4614 16438 4616 16490
rect 4616 16438 4668 16490
rect 4668 16438 4670 16490
rect 4614 16436 4670 16438
rect 4718 16490 4774 16492
rect 4718 16438 4720 16490
rect 4720 16438 4772 16490
rect 4772 16438 4774 16490
rect 4718 16436 4774 16438
rect 4822 16490 4878 16492
rect 4822 16438 4824 16490
rect 4824 16438 4876 16490
rect 4876 16438 4878 16490
rect 4822 16436 4878 16438
rect 11418 16490 11474 16492
rect 11418 16438 11420 16490
rect 11420 16438 11472 16490
rect 11472 16438 11474 16490
rect 11418 16436 11474 16438
rect 11522 16490 11578 16492
rect 11522 16438 11524 16490
rect 11524 16438 11576 16490
rect 11576 16438 11578 16490
rect 11522 16436 11578 16438
rect 11626 16490 11682 16492
rect 11626 16438 11628 16490
rect 11628 16438 11680 16490
rect 11680 16438 11682 16490
rect 11626 16436 11682 16438
rect 7196 16210 7252 16212
rect 7196 16158 7198 16210
rect 7198 16158 7250 16210
rect 7250 16158 7252 16210
rect 7196 16156 7252 16158
rect 10444 16156 10500 16212
rect 4956 15932 5012 15988
rect 5852 15986 5908 15988
rect 5852 15934 5854 15986
rect 5854 15934 5906 15986
rect 5906 15934 5908 15986
rect 5852 15932 5908 15934
rect 8016 15706 8072 15708
rect 8016 15654 8018 15706
rect 8018 15654 8070 15706
rect 8070 15654 8072 15706
rect 8016 15652 8072 15654
rect 8120 15706 8176 15708
rect 8120 15654 8122 15706
rect 8122 15654 8174 15706
rect 8174 15654 8176 15706
rect 8120 15652 8176 15654
rect 8224 15706 8280 15708
rect 8224 15654 8226 15706
rect 8226 15654 8278 15706
rect 8278 15654 8280 15706
rect 8224 15652 8280 15654
rect 4614 14922 4670 14924
rect 4614 14870 4616 14922
rect 4616 14870 4668 14922
rect 4668 14870 4670 14922
rect 4614 14868 4670 14870
rect 4718 14922 4774 14924
rect 4718 14870 4720 14922
rect 4720 14870 4772 14922
rect 4772 14870 4774 14922
rect 4718 14868 4774 14870
rect 4822 14922 4878 14924
rect 4822 14870 4824 14922
rect 4824 14870 4876 14922
rect 4876 14870 4878 14922
rect 4822 14868 4878 14870
rect 8016 14138 8072 14140
rect 8016 14086 8018 14138
rect 8018 14086 8070 14138
rect 8070 14086 8072 14138
rect 8016 14084 8072 14086
rect 8120 14138 8176 14140
rect 8120 14086 8122 14138
rect 8122 14086 8174 14138
rect 8174 14086 8176 14138
rect 8120 14084 8176 14086
rect 8224 14138 8280 14140
rect 8224 14086 8226 14138
rect 8226 14086 8278 14138
rect 8278 14086 8280 14138
rect 8224 14084 8280 14086
rect 4614 13354 4670 13356
rect 4614 13302 4616 13354
rect 4616 13302 4668 13354
rect 4668 13302 4670 13354
rect 4614 13300 4670 13302
rect 4718 13354 4774 13356
rect 4718 13302 4720 13354
rect 4720 13302 4772 13354
rect 4772 13302 4774 13354
rect 4718 13300 4774 13302
rect 4822 13354 4878 13356
rect 4822 13302 4824 13354
rect 4824 13302 4876 13354
rect 4876 13302 4878 13354
rect 4822 13300 4878 13302
rect 1708 12178 1764 12180
rect 1708 12126 1710 12178
rect 1710 12126 1762 12178
rect 1762 12126 1764 12178
rect 1708 12124 1764 12126
rect 7084 12850 7140 12852
rect 7084 12798 7086 12850
rect 7086 12798 7138 12850
rect 7138 12798 7140 12850
rect 7084 12796 7140 12798
rect 7644 12850 7700 12852
rect 7644 12798 7646 12850
rect 7646 12798 7698 12850
rect 7698 12798 7700 12850
rect 7644 12796 7700 12798
rect 7196 12738 7252 12740
rect 7196 12686 7198 12738
rect 7198 12686 7250 12738
rect 7250 12686 7252 12738
rect 7196 12684 7252 12686
rect 8016 12570 8072 12572
rect 8016 12518 8018 12570
rect 8018 12518 8070 12570
rect 8070 12518 8072 12570
rect 8016 12516 8072 12518
rect 8120 12570 8176 12572
rect 8120 12518 8122 12570
rect 8122 12518 8174 12570
rect 8174 12518 8176 12570
rect 8120 12516 8176 12518
rect 8224 12570 8280 12572
rect 8224 12518 8226 12570
rect 8226 12518 8278 12570
rect 8278 12518 8280 12570
rect 8224 12516 8280 12518
rect 3388 11900 3444 11956
rect 3612 11900 3668 11956
rect 3276 4562 3332 4564
rect 3276 4510 3278 4562
rect 3278 4510 3330 4562
rect 3330 4510 3332 4562
rect 3276 4508 3332 4510
rect 4614 11786 4670 11788
rect 4614 11734 4616 11786
rect 4616 11734 4668 11786
rect 4668 11734 4670 11786
rect 4614 11732 4670 11734
rect 4718 11786 4774 11788
rect 4718 11734 4720 11786
rect 4720 11734 4772 11786
rect 4772 11734 4774 11786
rect 4718 11732 4774 11734
rect 4822 11786 4878 11788
rect 4822 11734 4824 11786
rect 4824 11734 4876 11786
rect 4876 11734 4878 11786
rect 4822 11732 4878 11734
rect 8016 11002 8072 11004
rect 8016 10950 8018 11002
rect 8018 10950 8070 11002
rect 8070 10950 8072 11002
rect 8016 10948 8072 10950
rect 8120 11002 8176 11004
rect 8120 10950 8122 11002
rect 8122 10950 8174 11002
rect 8174 10950 8176 11002
rect 8120 10948 8176 10950
rect 8224 11002 8280 11004
rect 8224 10950 8226 11002
rect 8226 10950 8278 11002
rect 8278 10950 8280 11002
rect 8224 10948 8280 10950
rect 4614 10218 4670 10220
rect 4614 10166 4616 10218
rect 4616 10166 4668 10218
rect 4668 10166 4670 10218
rect 4614 10164 4670 10166
rect 4718 10218 4774 10220
rect 4718 10166 4720 10218
rect 4720 10166 4772 10218
rect 4772 10166 4774 10218
rect 4718 10164 4774 10166
rect 4822 10218 4878 10220
rect 4822 10166 4824 10218
rect 4824 10166 4876 10218
rect 4876 10166 4878 10218
rect 4822 10164 4878 10166
rect 8016 9434 8072 9436
rect 8016 9382 8018 9434
rect 8018 9382 8070 9434
rect 8070 9382 8072 9434
rect 8016 9380 8072 9382
rect 8120 9434 8176 9436
rect 8120 9382 8122 9434
rect 8122 9382 8174 9434
rect 8174 9382 8176 9434
rect 8120 9380 8176 9382
rect 8224 9434 8280 9436
rect 8224 9382 8226 9434
rect 8226 9382 8278 9434
rect 8278 9382 8280 9434
rect 8224 9380 8280 9382
rect 7756 8876 7812 8932
rect 4614 8650 4670 8652
rect 4614 8598 4616 8650
rect 4616 8598 4668 8650
rect 4668 8598 4670 8650
rect 4614 8596 4670 8598
rect 4718 8650 4774 8652
rect 4718 8598 4720 8650
rect 4720 8598 4772 8650
rect 4772 8598 4774 8650
rect 4718 8596 4774 8598
rect 4822 8650 4878 8652
rect 4822 8598 4824 8650
rect 4824 8598 4876 8650
rect 4876 8598 4878 8650
rect 4822 8596 4878 8598
rect 4614 7082 4670 7084
rect 4614 7030 4616 7082
rect 4616 7030 4668 7082
rect 4668 7030 4670 7082
rect 4614 7028 4670 7030
rect 4718 7082 4774 7084
rect 4718 7030 4720 7082
rect 4720 7030 4772 7082
rect 4772 7030 4774 7082
rect 4718 7028 4774 7030
rect 4822 7082 4878 7084
rect 4822 7030 4824 7082
rect 4824 7030 4876 7082
rect 4876 7030 4878 7082
rect 4822 7028 4878 7030
rect 7420 6860 7476 6916
rect 4614 5514 4670 5516
rect 4614 5462 4616 5514
rect 4616 5462 4668 5514
rect 4668 5462 4670 5514
rect 4614 5460 4670 5462
rect 4718 5514 4774 5516
rect 4718 5462 4720 5514
rect 4720 5462 4772 5514
rect 4772 5462 4774 5514
rect 4718 5460 4774 5462
rect 4822 5514 4878 5516
rect 4822 5462 4824 5514
rect 4824 5462 4876 5514
rect 4876 5462 4878 5514
rect 4822 5460 4878 5462
rect 6748 4844 6804 4900
rect 3612 4284 3668 4340
rect 4396 4396 4452 4452
rect 5180 4338 5236 4340
rect 5180 4286 5182 4338
rect 5182 4286 5234 4338
rect 5234 4286 5236 4338
rect 5180 4284 5236 4286
rect 5964 4338 6020 4340
rect 5964 4286 5966 4338
rect 5966 4286 6018 4338
rect 6018 4286 6020 4338
rect 5964 4284 6020 4286
rect 4614 3946 4670 3948
rect 4614 3894 4616 3946
rect 4616 3894 4668 3946
rect 4668 3894 4670 3946
rect 4614 3892 4670 3894
rect 4718 3946 4774 3948
rect 4718 3894 4720 3946
rect 4720 3894 4772 3946
rect 4772 3894 4774 3946
rect 4718 3892 4774 3894
rect 4822 3946 4878 3948
rect 4822 3894 4824 3946
rect 4824 3894 4876 3946
rect 4876 3894 4878 3946
rect 4822 3892 4878 3894
rect 7420 4508 7476 4564
rect 10108 8204 10164 8260
rect 8016 7866 8072 7868
rect 8016 7814 8018 7866
rect 8018 7814 8070 7866
rect 8070 7814 8072 7866
rect 8016 7812 8072 7814
rect 8120 7866 8176 7868
rect 8120 7814 8122 7866
rect 8122 7814 8174 7866
rect 8174 7814 8176 7866
rect 8120 7812 8176 7814
rect 8224 7866 8280 7868
rect 8224 7814 8226 7866
rect 8226 7814 8278 7866
rect 8278 7814 8280 7866
rect 8224 7812 8280 7814
rect 10108 6860 10164 6916
rect 16828 16210 16884 16212
rect 16828 16158 16830 16210
rect 16830 16158 16882 16210
rect 16882 16158 16884 16210
rect 16828 16156 16884 16158
rect 26460 17724 26516 17780
rect 18222 16490 18278 16492
rect 18222 16438 18224 16490
rect 18224 16438 18276 16490
rect 18276 16438 18278 16490
rect 18222 16436 18278 16438
rect 18326 16490 18382 16492
rect 18326 16438 18328 16490
rect 18328 16438 18380 16490
rect 18380 16438 18382 16490
rect 18326 16436 18382 16438
rect 18430 16490 18486 16492
rect 18430 16438 18432 16490
rect 18432 16438 18484 16490
rect 18484 16438 18486 16490
rect 18430 16436 18486 16438
rect 25026 16490 25082 16492
rect 25026 16438 25028 16490
rect 25028 16438 25080 16490
rect 25080 16438 25082 16490
rect 25026 16436 25082 16438
rect 25130 16490 25186 16492
rect 25130 16438 25132 16490
rect 25132 16438 25184 16490
rect 25184 16438 25186 16490
rect 25130 16436 25186 16438
rect 25234 16490 25290 16492
rect 25234 16438 25236 16490
rect 25236 16438 25288 16490
rect 25288 16438 25290 16490
rect 25234 16436 25290 16438
rect 17500 16156 17556 16212
rect 19740 16156 19796 16212
rect 29596 17724 29652 17780
rect 14820 15706 14876 15708
rect 14820 15654 14822 15706
rect 14822 15654 14874 15706
rect 14874 15654 14876 15706
rect 14820 15652 14876 15654
rect 14924 15706 14980 15708
rect 14924 15654 14926 15706
rect 14926 15654 14978 15706
rect 14978 15654 14980 15706
rect 14924 15652 14980 15654
rect 15028 15706 15084 15708
rect 15028 15654 15030 15706
rect 15030 15654 15082 15706
rect 15082 15654 15084 15706
rect 15028 15652 15084 15654
rect 14140 15484 14196 15540
rect 11418 14922 11474 14924
rect 11418 14870 11420 14922
rect 11420 14870 11472 14922
rect 11472 14870 11474 14922
rect 11418 14868 11474 14870
rect 11522 14922 11578 14924
rect 11522 14870 11524 14922
rect 11524 14870 11576 14922
rect 11576 14870 11578 14922
rect 11522 14868 11578 14870
rect 11626 14922 11682 14924
rect 11626 14870 11628 14922
rect 11628 14870 11680 14922
rect 11680 14870 11682 14922
rect 11626 14868 11682 14870
rect 14028 13468 14084 13524
rect 11418 13354 11474 13356
rect 11418 13302 11420 13354
rect 11420 13302 11472 13354
rect 11472 13302 11474 13354
rect 11418 13300 11474 13302
rect 11522 13354 11578 13356
rect 11522 13302 11524 13354
rect 11524 13302 11576 13354
rect 11576 13302 11578 13354
rect 11522 13300 11578 13302
rect 11626 13354 11682 13356
rect 11626 13302 11628 13354
rect 11628 13302 11680 13354
rect 11680 13302 11682 13354
rect 11626 13300 11682 13302
rect 13580 12684 13636 12740
rect 12796 11900 12852 11956
rect 11418 11786 11474 11788
rect 11418 11734 11420 11786
rect 11420 11734 11472 11786
rect 11472 11734 11474 11786
rect 11418 11732 11474 11734
rect 11522 11786 11578 11788
rect 11522 11734 11524 11786
rect 11524 11734 11576 11786
rect 11576 11734 11578 11786
rect 11522 11732 11578 11734
rect 11626 11786 11682 11788
rect 11626 11734 11628 11786
rect 11628 11734 11680 11786
rect 11680 11734 11682 11786
rect 11626 11732 11682 11734
rect 14820 14138 14876 14140
rect 14820 14086 14822 14138
rect 14822 14086 14874 14138
rect 14874 14086 14876 14138
rect 14820 14084 14876 14086
rect 14924 14138 14980 14140
rect 14924 14086 14926 14138
rect 14926 14086 14978 14138
rect 14978 14086 14980 14138
rect 14924 14084 14980 14086
rect 15028 14138 15084 14140
rect 15028 14086 15030 14138
rect 15030 14086 15082 14138
rect 15082 14086 15084 14138
rect 15028 14084 15084 14086
rect 21624 15706 21680 15708
rect 21624 15654 21626 15706
rect 21626 15654 21678 15706
rect 21678 15654 21680 15706
rect 21624 15652 21680 15654
rect 21728 15706 21784 15708
rect 21728 15654 21730 15706
rect 21730 15654 21782 15706
rect 21782 15654 21784 15706
rect 21728 15652 21784 15654
rect 21832 15706 21888 15708
rect 21832 15654 21834 15706
rect 21834 15654 21886 15706
rect 21886 15654 21888 15706
rect 21832 15652 21888 15654
rect 24556 15484 24612 15540
rect 28428 15706 28484 15708
rect 28428 15654 28430 15706
rect 28430 15654 28482 15706
rect 28482 15654 28484 15706
rect 28428 15652 28484 15654
rect 28532 15706 28588 15708
rect 28532 15654 28534 15706
rect 28534 15654 28586 15706
rect 28586 15654 28588 15706
rect 28532 15652 28588 15654
rect 28636 15706 28692 15708
rect 28636 15654 28638 15706
rect 28638 15654 28690 15706
rect 28690 15654 28692 15706
rect 28636 15652 28692 15654
rect 25340 15484 25396 15540
rect 18222 14922 18278 14924
rect 18222 14870 18224 14922
rect 18224 14870 18276 14922
rect 18276 14870 18278 14922
rect 18222 14868 18278 14870
rect 18326 14922 18382 14924
rect 18326 14870 18328 14922
rect 18328 14870 18380 14922
rect 18380 14870 18382 14922
rect 18326 14868 18382 14870
rect 18430 14922 18486 14924
rect 18430 14870 18432 14922
rect 18432 14870 18484 14922
rect 18484 14870 18486 14922
rect 18430 14868 18486 14870
rect 25026 14922 25082 14924
rect 25026 14870 25028 14922
rect 25028 14870 25080 14922
rect 25080 14870 25082 14922
rect 25026 14868 25082 14870
rect 25130 14922 25186 14924
rect 25130 14870 25132 14922
rect 25132 14870 25184 14922
rect 25184 14870 25186 14922
rect 25130 14868 25186 14870
rect 25234 14922 25290 14924
rect 25234 14870 25236 14922
rect 25236 14870 25288 14922
rect 25288 14870 25290 14922
rect 25234 14868 25290 14870
rect 21624 14138 21680 14140
rect 21624 14086 21626 14138
rect 21626 14086 21678 14138
rect 21678 14086 21680 14138
rect 21624 14084 21680 14086
rect 21728 14138 21784 14140
rect 21728 14086 21730 14138
rect 21730 14086 21782 14138
rect 21782 14086 21784 14138
rect 21728 14084 21784 14086
rect 21832 14138 21888 14140
rect 21832 14086 21834 14138
rect 21834 14086 21886 14138
rect 21886 14086 21888 14138
rect 21832 14084 21888 14086
rect 28428 14138 28484 14140
rect 28428 14086 28430 14138
rect 28430 14086 28482 14138
rect 28482 14086 28484 14138
rect 28428 14084 28484 14086
rect 28532 14138 28588 14140
rect 28532 14086 28534 14138
rect 28534 14086 28586 14138
rect 28586 14086 28588 14138
rect 28532 14084 28588 14086
rect 28636 14138 28692 14140
rect 28636 14086 28638 14138
rect 28638 14086 28690 14138
rect 28690 14086 28692 14138
rect 28636 14084 28692 14086
rect 15708 13804 15764 13860
rect 10556 8930 10612 8932
rect 10556 8878 10558 8930
rect 10558 8878 10610 8930
rect 10610 8878 10612 8930
rect 10556 8876 10612 8878
rect 14476 12796 14532 12852
rect 14820 12570 14876 12572
rect 14820 12518 14822 12570
rect 14822 12518 14874 12570
rect 14874 12518 14876 12570
rect 14820 12516 14876 12518
rect 14924 12570 14980 12572
rect 14924 12518 14926 12570
rect 14926 12518 14978 12570
rect 14978 12518 14980 12570
rect 14924 12516 14980 12518
rect 15028 12570 15084 12572
rect 15028 12518 15030 12570
rect 15030 12518 15082 12570
rect 15082 12518 15084 12570
rect 15028 12516 15084 12518
rect 10556 8428 10612 8484
rect 13100 8459 13156 8484
rect 13100 8428 13102 8459
rect 13102 8428 13154 8459
rect 13154 8428 13156 8459
rect 13100 8244 13102 8260
rect 13102 8244 13154 8260
rect 13154 8244 13156 8260
rect 13100 8204 13156 8244
rect 10444 8092 10500 8148
rect 12796 8121 12852 8148
rect 12796 8092 12798 8121
rect 12798 8092 12850 8121
rect 12850 8092 12852 8121
rect 8016 6298 8072 6300
rect 8016 6246 8018 6298
rect 8018 6246 8070 6298
rect 8070 6246 8072 6298
rect 8016 6244 8072 6246
rect 8120 6298 8176 6300
rect 8120 6246 8122 6298
rect 8122 6246 8174 6298
rect 8174 6246 8176 6298
rect 8120 6244 8176 6246
rect 8224 6298 8280 6300
rect 8224 6246 8226 6298
rect 8226 6246 8278 6298
rect 8278 6246 8280 6298
rect 8224 6244 8280 6246
rect 7868 4844 7924 4900
rect 15260 11900 15316 11956
rect 14820 11002 14876 11004
rect 14820 10950 14822 11002
rect 14822 10950 14874 11002
rect 14874 10950 14876 11002
rect 14820 10948 14876 10950
rect 14924 11002 14980 11004
rect 14924 10950 14926 11002
rect 14926 10950 14978 11002
rect 14978 10950 14980 11002
rect 14924 10948 14980 10950
rect 15028 11002 15084 11004
rect 15028 10950 15030 11002
rect 15030 10950 15082 11002
rect 15082 10950 15084 11002
rect 15028 10948 15084 10950
rect 14924 8121 14980 8148
rect 14924 8092 14926 8121
rect 14926 8092 14978 8121
rect 14978 8092 14980 8121
rect 11418 5514 11474 5516
rect 11418 5462 11420 5514
rect 11420 5462 11472 5514
rect 11472 5462 11474 5514
rect 11418 5460 11474 5462
rect 11522 5514 11578 5516
rect 11522 5462 11524 5514
rect 11524 5462 11576 5514
rect 11576 5462 11578 5514
rect 11522 5460 11578 5462
rect 11626 5514 11682 5516
rect 11626 5462 11628 5514
rect 11628 5462 11680 5514
rect 11680 5462 11682 5514
rect 11626 5460 11682 5462
rect 10444 4844 10500 4900
rect 8016 4730 8072 4732
rect 8016 4678 8018 4730
rect 8018 4678 8070 4730
rect 8070 4678 8072 4730
rect 8016 4676 8072 4678
rect 8120 4730 8176 4732
rect 8120 4678 8122 4730
rect 8122 4678 8174 4730
rect 8174 4678 8176 4730
rect 8120 4676 8176 4678
rect 8224 4730 8280 4732
rect 8224 4678 8226 4730
rect 8226 4678 8278 4730
rect 8278 4678 8280 4730
rect 8224 4676 8280 4678
rect 8764 4562 8820 4564
rect 8764 4510 8766 4562
rect 8766 4510 8818 4562
rect 8818 4510 8820 4562
rect 8764 4508 8820 4510
rect 7756 4396 7812 4452
rect 7084 4172 7140 4228
rect 8316 4338 8372 4340
rect 8316 4286 8318 4338
rect 8318 4286 8370 4338
rect 8370 4286 8372 4338
rect 8316 4284 8372 4286
rect 8764 4172 8820 4228
rect 14820 4730 14876 4732
rect 14820 4678 14822 4730
rect 14822 4678 14874 4730
rect 14874 4678 14876 4730
rect 14820 4676 14876 4678
rect 14924 4730 14980 4732
rect 14924 4678 14926 4730
rect 14926 4678 14978 4730
rect 14978 4678 14980 4730
rect 14924 4676 14980 4678
rect 15028 4730 15084 4732
rect 15028 4678 15030 4730
rect 15030 4678 15082 4730
rect 15082 4678 15084 4730
rect 15028 4676 15084 4678
rect 16604 13858 16660 13860
rect 16604 13806 16606 13858
rect 16606 13806 16658 13858
rect 16658 13806 16660 13858
rect 16604 13804 16660 13806
rect 17612 13804 17668 13860
rect 16492 13522 16548 13524
rect 16492 13470 16494 13522
rect 16494 13470 16546 13522
rect 16546 13470 16548 13522
rect 16492 13468 16548 13470
rect 18222 13354 18278 13356
rect 18222 13302 18224 13354
rect 18224 13302 18276 13354
rect 18276 13302 18278 13354
rect 18222 13300 18278 13302
rect 18326 13354 18382 13356
rect 18326 13302 18328 13354
rect 18328 13302 18380 13354
rect 18380 13302 18382 13354
rect 18326 13300 18382 13302
rect 18430 13354 18486 13356
rect 18430 13302 18432 13354
rect 18432 13302 18484 13354
rect 18484 13302 18486 13354
rect 18430 13300 18486 13302
rect 25026 13354 25082 13356
rect 25026 13302 25028 13354
rect 25028 13302 25080 13354
rect 25080 13302 25082 13354
rect 25026 13300 25082 13302
rect 25130 13354 25186 13356
rect 25130 13302 25132 13354
rect 25132 13302 25184 13354
rect 25184 13302 25186 13354
rect 25130 13300 25186 13302
rect 25234 13354 25290 13356
rect 25234 13302 25236 13354
rect 25236 13302 25288 13354
rect 25288 13302 25290 13354
rect 25234 13300 25290 13302
rect 21624 12570 21680 12572
rect 21624 12518 21626 12570
rect 21626 12518 21678 12570
rect 21678 12518 21680 12570
rect 21624 12516 21680 12518
rect 21728 12570 21784 12572
rect 21728 12518 21730 12570
rect 21730 12518 21782 12570
rect 21782 12518 21784 12570
rect 21728 12516 21784 12518
rect 21832 12570 21888 12572
rect 21832 12518 21834 12570
rect 21834 12518 21886 12570
rect 21886 12518 21888 12570
rect 21832 12516 21888 12518
rect 28428 12570 28484 12572
rect 28428 12518 28430 12570
rect 28430 12518 28482 12570
rect 28482 12518 28484 12570
rect 28428 12516 28484 12518
rect 28532 12570 28588 12572
rect 28532 12518 28534 12570
rect 28534 12518 28586 12570
rect 28586 12518 28588 12570
rect 28532 12516 28588 12518
rect 28636 12570 28692 12572
rect 28636 12518 28638 12570
rect 28638 12518 28690 12570
rect 28690 12518 28692 12570
rect 28636 12516 28692 12518
rect 18222 11786 18278 11788
rect 18222 11734 18224 11786
rect 18224 11734 18276 11786
rect 18276 11734 18278 11786
rect 18222 11732 18278 11734
rect 18326 11786 18382 11788
rect 18326 11734 18328 11786
rect 18328 11734 18380 11786
rect 18380 11734 18382 11786
rect 18326 11732 18382 11734
rect 18430 11786 18486 11788
rect 18430 11734 18432 11786
rect 18432 11734 18484 11786
rect 18484 11734 18486 11786
rect 18430 11732 18486 11734
rect 25026 11786 25082 11788
rect 25026 11734 25028 11786
rect 25028 11734 25080 11786
rect 25080 11734 25082 11786
rect 25026 11732 25082 11734
rect 25130 11786 25186 11788
rect 25130 11734 25132 11786
rect 25132 11734 25184 11786
rect 25184 11734 25186 11786
rect 25130 11732 25186 11734
rect 25234 11786 25290 11788
rect 25234 11734 25236 11786
rect 25236 11734 25288 11786
rect 25288 11734 25290 11786
rect 25234 11732 25290 11734
rect 21624 11002 21680 11004
rect 21624 10950 21626 11002
rect 21626 10950 21678 11002
rect 21678 10950 21680 11002
rect 21624 10948 21680 10950
rect 21728 11002 21784 11004
rect 21728 10950 21730 11002
rect 21730 10950 21782 11002
rect 21782 10950 21784 11002
rect 21728 10948 21784 10950
rect 21832 11002 21888 11004
rect 21832 10950 21834 11002
rect 21834 10950 21886 11002
rect 21886 10950 21888 11002
rect 21832 10948 21888 10950
rect 28428 11002 28484 11004
rect 28428 10950 28430 11002
rect 28430 10950 28482 11002
rect 28482 10950 28484 11002
rect 28428 10948 28484 10950
rect 28532 11002 28588 11004
rect 28532 10950 28534 11002
rect 28534 10950 28586 11002
rect 28586 10950 28588 11002
rect 28532 10948 28588 10950
rect 28636 11002 28692 11004
rect 28636 10950 28638 11002
rect 28638 10950 28690 11002
rect 28690 10950 28692 11002
rect 28636 10948 28692 10950
rect 18222 10218 18278 10220
rect 18222 10166 18224 10218
rect 18224 10166 18276 10218
rect 18276 10166 18278 10218
rect 18222 10164 18278 10166
rect 18326 10218 18382 10220
rect 18326 10166 18328 10218
rect 18328 10166 18380 10218
rect 18380 10166 18382 10218
rect 18326 10164 18382 10166
rect 18430 10218 18486 10220
rect 18430 10166 18432 10218
rect 18432 10166 18484 10218
rect 18484 10166 18486 10218
rect 18430 10164 18486 10166
rect 25026 10218 25082 10220
rect 25026 10166 25028 10218
rect 25028 10166 25080 10218
rect 25080 10166 25082 10218
rect 25026 10164 25082 10166
rect 25130 10218 25186 10220
rect 25130 10166 25132 10218
rect 25132 10166 25184 10218
rect 25184 10166 25186 10218
rect 25130 10164 25186 10166
rect 25234 10218 25290 10220
rect 25234 10166 25236 10218
rect 25236 10166 25288 10218
rect 25288 10166 25290 10218
rect 25234 10164 25290 10166
rect 21624 9434 21680 9436
rect 21624 9382 21626 9434
rect 21626 9382 21678 9434
rect 21678 9382 21680 9434
rect 21624 9380 21680 9382
rect 21728 9434 21784 9436
rect 21728 9382 21730 9434
rect 21730 9382 21782 9434
rect 21782 9382 21784 9434
rect 21728 9380 21784 9382
rect 21832 9434 21888 9436
rect 21832 9382 21834 9434
rect 21834 9382 21886 9434
rect 21886 9382 21888 9434
rect 21832 9380 21888 9382
rect 28428 9434 28484 9436
rect 28428 9382 28430 9434
rect 28430 9382 28482 9434
rect 28482 9382 28484 9434
rect 28428 9380 28484 9382
rect 28532 9434 28588 9436
rect 28532 9382 28534 9434
rect 28534 9382 28586 9434
rect 28586 9382 28588 9434
rect 28532 9380 28588 9382
rect 28636 9434 28692 9436
rect 28636 9382 28638 9434
rect 28638 9382 28690 9434
rect 28690 9382 28692 9434
rect 28636 9380 28692 9382
rect 15462 8482 15518 8484
rect 15462 8430 15464 8482
rect 15464 8430 15516 8482
rect 15516 8430 15518 8482
rect 15462 8428 15518 8430
rect 18284 8764 18340 8820
rect 18222 8650 18278 8652
rect 18222 8598 18224 8650
rect 18224 8598 18276 8650
rect 18276 8598 18278 8650
rect 18222 8596 18278 8598
rect 18326 8650 18382 8652
rect 18326 8598 18328 8650
rect 18328 8598 18380 8650
rect 18380 8598 18382 8650
rect 18326 8596 18382 8598
rect 18430 8650 18486 8652
rect 18430 8598 18432 8650
rect 18432 8598 18484 8650
rect 18484 8598 18486 8650
rect 18430 8596 18486 8598
rect 18060 8428 18116 8484
rect 15467 8248 15469 8260
rect 15469 8248 15521 8260
rect 15521 8248 15523 8260
rect 15467 8204 15523 8248
rect 24892 8764 24948 8820
rect 25026 8650 25082 8652
rect 25026 8598 25028 8650
rect 25028 8598 25080 8650
rect 25080 8598 25082 8650
rect 25026 8596 25082 8598
rect 25130 8650 25186 8652
rect 25130 8598 25132 8650
rect 25132 8598 25184 8650
rect 25184 8598 25186 8650
rect 25130 8596 25186 8598
rect 25234 8650 25290 8652
rect 25234 8598 25236 8650
rect 25236 8598 25288 8650
rect 25288 8598 25290 8650
rect 25234 8596 25290 8598
rect 18620 8204 18676 8260
rect 18172 8146 18228 8148
rect 18172 8094 18174 8146
rect 18174 8094 18226 8146
rect 18226 8094 18228 8146
rect 18172 8092 18228 8094
rect 26236 8146 26292 8148
rect 26236 8094 26238 8146
rect 26238 8094 26290 8146
rect 26290 8094 26292 8146
rect 26236 8092 26292 8094
rect 26908 8092 26964 8148
rect 21624 7866 21680 7868
rect 21624 7814 21626 7866
rect 21626 7814 21678 7866
rect 21678 7814 21680 7866
rect 21624 7812 21680 7814
rect 21728 7866 21784 7868
rect 21728 7814 21730 7866
rect 21730 7814 21782 7866
rect 21782 7814 21784 7866
rect 21728 7812 21784 7814
rect 21832 7866 21888 7868
rect 21832 7814 21834 7866
rect 21834 7814 21886 7866
rect 21886 7814 21888 7866
rect 21832 7812 21888 7814
rect 28428 7866 28484 7868
rect 28428 7814 28430 7866
rect 28430 7814 28482 7866
rect 28482 7814 28484 7866
rect 28428 7812 28484 7814
rect 28532 7866 28588 7868
rect 28532 7814 28534 7866
rect 28534 7814 28586 7866
rect 28586 7814 28588 7866
rect 28532 7812 28588 7814
rect 28636 7866 28692 7868
rect 28636 7814 28638 7866
rect 28638 7814 28690 7866
rect 28690 7814 28692 7866
rect 28636 7812 28692 7814
rect 26908 7420 26964 7476
rect 18222 7082 18278 7084
rect 18222 7030 18224 7082
rect 18224 7030 18276 7082
rect 18276 7030 18278 7082
rect 18222 7028 18278 7030
rect 18326 7082 18382 7084
rect 18326 7030 18328 7082
rect 18328 7030 18380 7082
rect 18380 7030 18382 7082
rect 18326 7028 18382 7030
rect 18430 7082 18486 7084
rect 18430 7030 18432 7082
rect 18432 7030 18484 7082
rect 18484 7030 18486 7082
rect 18430 7028 18486 7030
rect 25026 7082 25082 7084
rect 25026 7030 25028 7082
rect 25028 7030 25080 7082
rect 25080 7030 25082 7082
rect 25026 7028 25082 7030
rect 25130 7082 25186 7084
rect 25130 7030 25132 7082
rect 25132 7030 25184 7082
rect 25184 7030 25186 7082
rect 25130 7028 25186 7030
rect 25234 7082 25290 7084
rect 25234 7030 25236 7082
rect 25236 7030 25288 7082
rect 25288 7030 25290 7082
rect 25234 7028 25290 7030
rect 21624 6298 21680 6300
rect 21624 6246 21626 6298
rect 21626 6246 21678 6298
rect 21678 6246 21680 6298
rect 21624 6244 21680 6246
rect 21728 6298 21784 6300
rect 21728 6246 21730 6298
rect 21730 6246 21782 6298
rect 21782 6246 21784 6298
rect 21728 6244 21784 6246
rect 21832 6298 21888 6300
rect 21832 6246 21834 6298
rect 21834 6246 21886 6298
rect 21886 6246 21888 6298
rect 21832 6244 21888 6246
rect 28428 6298 28484 6300
rect 28428 6246 28430 6298
rect 28430 6246 28482 6298
rect 28482 6246 28484 6298
rect 28428 6244 28484 6246
rect 28532 6298 28588 6300
rect 28532 6246 28534 6298
rect 28534 6246 28586 6298
rect 28586 6246 28588 6298
rect 28532 6244 28588 6246
rect 28636 6298 28692 6300
rect 28636 6246 28638 6298
rect 28638 6246 28690 6298
rect 28690 6246 28692 6298
rect 28636 6244 28692 6246
rect 18222 5514 18278 5516
rect 18222 5462 18224 5514
rect 18224 5462 18276 5514
rect 18276 5462 18278 5514
rect 18222 5460 18278 5462
rect 18326 5514 18382 5516
rect 18326 5462 18328 5514
rect 18328 5462 18380 5514
rect 18380 5462 18382 5514
rect 18326 5460 18382 5462
rect 18430 5514 18486 5516
rect 18430 5462 18432 5514
rect 18432 5462 18484 5514
rect 18484 5462 18486 5514
rect 18430 5460 18486 5462
rect 25026 5514 25082 5516
rect 25026 5462 25028 5514
rect 25028 5462 25080 5514
rect 25080 5462 25082 5514
rect 25026 5460 25082 5462
rect 25130 5514 25186 5516
rect 25130 5462 25132 5514
rect 25132 5462 25184 5514
rect 25184 5462 25186 5514
rect 25130 5460 25186 5462
rect 25234 5514 25290 5516
rect 25234 5462 25236 5514
rect 25236 5462 25288 5514
rect 25288 5462 25290 5514
rect 25234 5460 25290 5462
rect 21624 4730 21680 4732
rect 21624 4678 21626 4730
rect 21626 4678 21678 4730
rect 21678 4678 21680 4730
rect 21624 4676 21680 4678
rect 21728 4730 21784 4732
rect 21728 4678 21730 4730
rect 21730 4678 21782 4730
rect 21782 4678 21784 4730
rect 21728 4676 21784 4678
rect 21832 4730 21888 4732
rect 21832 4678 21834 4730
rect 21834 4678 21886 4730
rect 21886 4678 21888 4730
rect 21832 4676 21888 4678
rect 28428 4730 28484 4732
rect 28428 4678 28430 4730
rect 28430 4678 28482 4730
rect 28482 4678 28484 4730
rect 28428 4676 28484 4678
rect 28532 4730 28588 4732
rect 28532 4678 28534 4730
rect 28534 4678 28586 4730
rect 28586 4678 28588 4730
rect 28532 4676 28588 4678
rect 28636 4730 28692 4732
rect 28636 4678 28638 4730
rect 28638 4678 28690 4730
rect 28690 4678 28692 4730
rect 28636 4676 28692 4678
rect 15148 4508 15204 4564
rect 14476 4284 14532 4340
rect 11418 3946 11474 3948
rect 11418 3894 11420 3946
rect 11420 3894 11472 3946
rect 11472 3894 11474 3946
rect 11418 3892 11474 3894
rect 11522 3946 11578 3948
rect 11522 3894 11524 3946
rect 11524 3894 11576 3946
rect 11576 3894 11578 3946
rect 11522 3892 11578 3894
rect 11626 3946 11682 3948
rect 11626 3894 11628 3946
rect 11628 3894 11680 3946
rect 11680 3894 11682 3946
rect 11626 3892 11682 3894
rect 6412 3500 6468 3556
rect 11564 3554 11620 3556
rect 11564 3502 11566 3554
rect 11566 3502 11618 3554
rect 11618 3502 11620 3554
rect 11564 3500 11620 3502
rect 28 2492 84 2548
rect 8016 3162 8072 3164
rect 8016 3110 8018 3162
rect 8018 3110 8070 3162
rect 8070 3110 8072 3162
rect 8016 3108 8072 3110
rect 8120 3162 8176 3164
rect 8120 3110 8122 3162
rect 8122 3110 8174 3162
rect 8174 3110 8176 3162
rect 8120 3108 8176 3110
rect 8224 3162 8280 3164
rect 8224 3110 8226 3162
rect 8226 3110 8278 3162
rect 8278 3110 8280 3162
rect 8224 3108 8280 3110
rect 1932 2492 1988 2548
rect 18222 3946 18278 3948
rect 18222 3894 18224 3946
rect 18224 3894 18276 3946
rect 18276 3894 18278 3946
rect 18222 3892 18278 3894
rect 18326 3946 18382 3948
rect 18326 3894 18328 3946
rect 18328 3894 18380 3946
rect 18380 3894 18382 3946
rect 18326 3892 18382 3894
rect 18430 3946 18486 3948
rect 18430 3894 18432 3946
rect 18432 3894 18484 3946
rect 18484 3894 18486 3946
rect 18430 3892 18486 3894
rect 25026 3946 25082 3948
rect 25026 3894 25028 3946
rect 25028 3894 25080 3946
rect 25080 3894 25082 3946
rect 25026 3892 25082 3894
rect 25130 3946 25186 3948
rect 25130 3894 25132 3946
rect 25132 3894 25184 3946
rect 25184 3894 25186 3946
rect 25130 3892 25186 3894
rect 25234 3946 25290 3948
rect 25234 3894 25236 3946
rect 25236 3894 25288 3946
rect 25288 3894 25290 3946
rect 25234 3892 25290 3894
rect 14476 3612 14532 3668
rect 25340 3666 25396 3668
rect 25340 3614 25342 3666
rect 25342 3614 25394 3666
rect 25394 3614 25396 3666
rect 25340 3612 25396 3614
rect 24892 3388 24948 3444
rect 14820 3162 14876 3164
rect 14820 3110 14822 3162
rect 14822 3110 14874 3162
rect 14874 3110 14876 3162
rect 14820 3108 14876 3110
rect 14924 3162 14980 3164
rect 14924 3110 14926 3162
rect 14926 3110 14978 3162
rect 14978 3110 14980 3162
rect 14924 3108 14980 3110
rect 15028 3162 15084 3164
rect 15028 3110 15030 3162
rect 15030 3110 15082 3162
rect 15082 3110 15084 3162
rect 15028 3108 15084 3110
rect 21624 3162 21680 3164
rect 21624 3110 21626 3162
rect 21626 3110 21678 3162
rect 21678 3110 21680 3162
rect 21624 3108 21680 3110
rect 21728 3162 21784 3164
rect 21728 3110 21730 3162
rect 21730 3110 21782 3162
rect 21782 3110 21784 3162
rect 21728 3108 21784 3110
rect 21832 3162 21888 3164
rect 21832 3110 21834 3162
rect 21834 3110 21886 3162
rect 21886 3110 21888 3162
rect 21832 3108 21888 3110
rect 26348 3442 26404 3444
rect 26348 3390 26350 3442
rect 26350 3390 26402 3442
rect 26402 3390 26404 3442
rect 26348 3388 26404 3390
rect 28428 3162 28484 3164
rect 28428 3110 28430 3162
rect 28430 3110 28482 3162
rect 28482 3110 28484 3162
rect 28428 3108 28484 3110
rect 28532 3162 28588 3164
rect 28532 3110 28534 3162
rect 28534 3110 28586 3162
rect 28586 3110 28588 3162
rect 28532 3108 28588 3110
rect 28636 3162 28692 3164
rect 28636 3110 28638 3162
rect 28638 3110 28690 3162
rect 28690 3110 28692 3162
rect 28636 3108 28692 3110
<< metal3 >>
rect 26450 17724 26460 17780
rect 26516 17724 29596 17780
rect 29652 17724 29662 17780
rect 4604 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4888 16492
rect 11408 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11692 16492
rect 18212 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18496 16492
rect 25016 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25300 16492
rect 7186 16156 7196 16212
rect 7252 16156 10444 16212
rect 10500 16156 10510 16212
rect 16818 16156 16828 16212
rect 16884 16156 17500 16212
rect 17556 16156 19740 16212
rect 19796 16156 19806 16212
rect 4946 15932 4956 15988
rect 5012 15932 5852 15988
rect 5908 15932 5918 15988
rect 8006 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8290 15708
rect 14810 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15094 15708
rect 21614 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21898 15708
rect 28418 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28702 15708
rect 14130 15484 14140 15540
rect 14196 15484 24556 15540
rect 24612 15484 25340 15540
rect 25396 15484 25406 15540
rect 4604 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4888 14924
rect 11408 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11692 14924
rect 18212 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18496 14924
rect 25016 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25300 14924
rect 8006 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8290 14140
rect 14810 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15094 14140
rect 21614 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21898 14140
rect 28418 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28702 14140
rect 15698 13804 15708 13860
rect 15764 13804 16604 13860
rect 16660 13804 17612 13860
rect 17668 13804 17678 13860
rect 14018 13468 14028 13524
rect 14084 13468 16492 13524
rect 16548 13468 16558 13524
rect 4604 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4888 13356
rect 11408 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11692 13356
rect 18212 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18496 13356
rect 25016 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25300 13356
rect 7074 12796 7084 12852
rect 7140 12796 7644 12852
rect 7700 12796 14476 12852
rect 14532 12796 14542 12852
rect 7186 12684 7196 12740
rect 7252 12684 13580 12740
rect 13636 12684 13646 12740
rect 8006 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8290 12572
rect 14810 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15094 12572
rect 21614 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21898 12572
rect 28418 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28702 12572
rect 200 12180 800 12208
rect 200 12124 1708 12180
rect 1764 12124 1774 12180
rect 200 12096 800 12124
rect 3378 11900 3388 11956
rect 3444 11900 3612 11956
rect 3668 11900 12796 11956
rect 12852 11900 15260 11956
rect 15316 11900 15326 11956
rect 4604 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4888 11788
rect 11408 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11692 11788
rect 18212 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18496 11788
rect 25016 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25300 11788
rect 8006 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8290 11004
rect 14810 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15094 11004
rect 21614 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21898 11004
rect 28418 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28702 11004
rect 4604 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4888 10220
rect 18212 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18496 10220
rect 25016 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25300 10220
rect 8006 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8290 9436
rect 21614 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21898 9436
rect 28418 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28702 9436
rect 7746 8876 7756 8932
rect 7812 8876 10556 8932
rect 10612 8876 10622 8932
rect 18274 8764 18284 8820
rect 18340 8764 24892 8820
rect 24948 8764 24958 8820
rect 4604 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4888 8652
rect 18212 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18496 8652
rect 25016 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25300 8652
rect 10546 8428 10556 8484
rect 10612 8428 13100 8484
rect 13156 8428 15462 8484
rect 15518 8428 18060 8484
rect 18116 8428 18126 8484
rect 10098 8204 10108 8260
rect 10164 8204 13100 8260
rect 13156 8204 15467 8260
rect 15523 8204 18620 8260
rect 18676 8204 18686 8260
rect 10434 8092 10444 8148
rect 10500 8092 12796 8148
rect 12852 8092 14924 8148
rect 14980 8092 18172 8148
rect 18228 8092 18238 8148
rect 26226 8092 26236 8148
rect 26292 8092 26908 8148
rect 26964 8092 26974 8148
rect 8006 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8290 7868
rect 21614 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21898 7868
rect 28418 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28702 7868
rect 29200 7476 29800 7504
rect 26898 7420 26908 7476
rect 26964 7420 29800 7476
rect 29200 7392 29800 7420
rect 4604 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4888 7084
rect 18212 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18496 7084
rect 25016 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25300 7084
rect 7410 6860 7420 6916
rect 7476 6860 10108 6916
rect 10164 6860 10174 6916
rect 8006 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8290 6300
rect 21614 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21898 6300
rect 28418 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28702 6300
rect 4604 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4888 5516
rect 11408 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11692 5516
rect 18212 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18496 5516
rect 25016 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25300 5516
rect 6738 4844 6748 4900
rect 6804 4844 7868 4900
rect 7924 4844 10444 4900
rect 10500 4844 10510 4900
rect 8006 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8290 4732
rect 14810 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15094 4732
rect 21614 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21898 4732
rect 28418 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28702 4732
rect 3266 4508 3276 4564
rect 3332 4508 7420 4564
rect 7476 4508 7486 4564
rect 8754 4508 8764 4564
rect 8820 4508 15148 4564
rect 15204 4508 15214 4564
rect 4386 4396 4396 4452
rect 4452 4396 7756 4452
rect 7812 4396 7822 4452
rect 3602 4284 3612 4340
rect 3668 4284 5180 4340
rect 5236 4284 5246 4340
rect 5954 4284 5964 4340
rect 6020 4284 8316 4340
rect 8372 4284 14476 4340
rect 14532 4284 14542 4340
rect 7074 4172 7084 4228
rect 7140 4172 8764 4228
rect 8820 4172 8830 4228
rect 4604 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4888 3948
rect 11408 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11692 3948
rect 18212 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18496 3948
rect 25016 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25300 3948
rect 14466 3612 14476 3668
rect 14532 3612 25340 3668
rect 25396 3612 25406 3668
rect 6402 3500 6412 3556
rect 6468 3500 11564 3556
rect 11620 3500 11630 3556
rect 24882 3388 24892 3444
rect 24948 3388 26348 3444
rect 26404 3388 26414 3444
rect 8006 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8290 3164
rect 14810 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15094 3164
rect 21614 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21898 3164
rect 28418 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28702 3164
rect 18 2492 28 2548
rect 84 2492 1932 2548
rect 1988 2492 1998 2548
<< via3 >>
rect 4614 16436 4670 16492
rect 4718 16436 4774 16492
rect 4822 16436 4878 16492
rect 11418 16436 11474 16492
rect 11522 16436 11578 16492
rect 11626 16436 11682 16492
rect 18222 16436 18278 16492
rect 18326 16436 18382 16492
rect 18430 16436 18486 16492
rect 25026 16436 25082 16492
rect 25130 16436 25186 16492
rect 25234 16436 25290 16492
rect 8016 15652 8072 15708
rect 8120 15652 8176 15708
rect 8224 15652 8280 15708
rect 14820 15652 14876 15708
rect 14924 15652 14980 15708
rect 15028 15652 15084 15708
rect 21624 15652 21680 15708
rect 21728 15652 21784 15708
rect 21832 15652 21888 15708
rect 28428 15652 28484 15708
rect 28532 15652 28588 15708
rect 28636 15652 28692 15708
rect 4614 14868 4670 14924
rect 4718 14868 4774 14924
rect 4822 14868 4878 14924
rect 11418 14868 11474 14924
rect 11522 14868 11578 14924
rect 11626 14868 11682 14924
rect 18222 14868 18278 14924
rect 18326 14868 18382 14924
rect 18430 14868 18486 14924
rect 25026 14868 25082 14924
rect 25130 14868 25186 14924
rect 25234 14868 25290 14924
rect 8016 14084 8072 14140
rect 8120 14084 8176 14140
rect 8224 14084 8280 14140
rect 14820 14084 14876 14140
rect 14924 14084 14980 14140
rect 15028 14084 15084 14140
rect 21624 14084 21680 14140
rect 21728 14084 21784 14140
rect 21832 14084 21888 14140
rect 28428 14084 28484 14140
rect 28532 14084 28588 14140
rect 28636 14084 28692 14140
rect 4614 13300 4670 13356
rect 4718 13300 4774 13356
rect 4822 13300 4878 13356
rect 11418 13300 11474 13356
rect 11522 13300 11578 13356
rect 11626 13300 11682 13356
rect 18222 13300 18278 13356
rect 18326 13300 18382 13356
rect 18430 13300 18486 13356
rect 25026 13300 25082 13356
rect 25130 13300 25186 13356
rect 25234 13300 25290 13356
rect 8016 12516 8072 12572
rect 8120 12516 8176 12572
rect 8224 12516 8280 12572
rect 14820 12516 14876 12572
rect 14924 12516 14980 12572
rect 15028 12516 15084 12572
rect 21624 12516 21680 12572
rect 21728 12516 21784 12572
rect 21832 12516 21888 12572
rect 28428 12516 28484 12572
rect 28532 12516 28588 12572
rect 28636 12516 28692 12572
rect 4614 11732 4670 11788
rect 4718 11732 4774 11788
rect 4822 11732 4878 11788
rect 11418 11732 11474 11788
rect 11522 11732 11578 11788
rect 11626 11732 11682 11788
rect 18222 11732 18278 11788
rect 18326 11732 18382 11788
rect 18430 11732 18486 11788
rect 25026 11732 25082 11788
rect 25130 11732 25186 11788
rect 25234 11732 25290 11788
rect 8016 10948 8072 11004
rect 8120 10948 8176 11004
rect 8224 10948 8280 11004
rect 14820 10948 14876 11004
rect 14924 10948 14980 11004
rect 15028 10948 15084 11004
rect 21624 10948 21680 11004
rect 21728 10948 21784 11004
rect 21832 10948 21888 11004
rect 28428 10948 28484 11004
rect 28532 10948 28588 11004
rect 28636 10948 28692 11004
rect 4614 10164 4670 10220
rect 4718 10164 4774 10220
rect 4822 10164 4878 10220
rect 18222 10164 18278 10220
rect 18326 10164 18382 10220
rect 18430 10164 18486 10220
rect 25026 10164 25082 10220
rect 25130 10164 25186 10220
rect 25234 10164 25290 10220
rect 8016 9380 8072 9436
rect 8120 9380 8176 9436
rect 8224 9380 8280 9436
rect 21624 9380 21680 9436
rect 21728 9380 21784 9436
rect 21832 9380 21888 9436
rect 28428 9380 28484 9436
rect 28532 9380 28588 9436
rect 28636 9380 28692 9436
rect 4614 8596 4670 8652
rect 4718 8596 4774 8652
rect 4822 8596 4878 8652
rect 18222 8596 18278 8652
rect 18326 8596 18382 8652
rect 18430 8596 18486 8652
rect 25026 8596 25082 8652
rect 25130 8596 25186 8652
rect 25234 8596 25290 8652
rect 8016 7812 8072 7868
rect 8120 7812 8176 7868
rect 8224 7812 8280 7868
rect 21624 7812 21680 7868
rect 21728 7812 21784 7868
rect 21832 7812 21888 7868
rect 28428 7812 28484 7868
rect 28532 7812 28588 7868
rect 28636 7812 28692 7868
rect 4614 7028 4670 7084
rect 4718 7028 4774 7084
rect 4822 7028 4878 7084
rect 18222 7028 18278 7084
rect 18326 7028 18382 7084
rect 18430 7028 18486 7084
rect 25026 7028 25082 7084
rect 25130 7028 25186 7084
rect 25234 7028 25290 7084
rect 8016 6244 8072 6300
rect 8120 6244 8176 6300
rect 8224 6244 8280 6300
rect 21624 6244 21680 6300
rect 21728 6244 21784 6300
rect 21832 6244 21888 6300
rect 28428 6244 28484 6300
rect 28532 6244 28588 6300
rect 28636 6244 28692 6300
rect 4614 5460 4670 5516
rect 4718 5460 4774 5516
rect 4822 5460 4878 5516
rect 11418 5460 11474 5516
rect 11522 5460 11578 5516
rect 11626 5460 11682 5516
rect 18222 5460 18278 5516
rect 18326 5460 18382 5516
rect 18430 5460 18486 5516
rect 25026 5460 25082 5516
rect 25130 5460 25186 5516
rect 25234 5460 25290 5516
rect 8016 4676 8072 4732
rect 8120 4676 8176 4732
rect 8224 4676 8280 4732
rect 14820 4676 14876 4732
rect 14924 4676 14980 4732
rect 15028 4676 15084 4732
rect 21624 4676 21680 4732
rect 21728 4676 21784 4732
rect 21832 4676 21888 4732
rect 28428 4676 28484 4732
rect 28532 4676 28588 4732
rect 28636 4676 28692 4732
rect 4614 3892 4670 3948
rect 4718 3892 4774 3948
rect 4822 3892 4878 3948
rect 11418 3892 11474 3948
rect 11522 3892 11578 3948
rect 11626 3892 11682 3948
rect 18222 3892 18278 3948
rect 18326 3892 18382 3948
rect 18430 3892 18486 3948
rect 25026 3892 25082 3948
rect 25130 3892 25186 3948
rect 25234 3892 25290 3948
rect 8016 3108 8072 3164
rect 8120 3108 8176 3164
rect 8224 3108 8280 3164
rect 14820 3108 14876 3164
rect 14924 3108 14980 3164
rect 15028 3108 15084 3164
rect 21624 3108 21680 3164
rect 21728 3108 21784 3164
rect 21832 3108 21888 3164
rect 28428 3108 28484 3164
rect 28532 3108 28588 3164
rect 28636 3108 28692 3164
<< metal4 >>
rect 4586 16492 4906 16524
rect 4586 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4906 16492
rect 4586 14924 4906 16436
rect 4586 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4906 14924
rect 4586 13356 4906 14868
rect 4586 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4906 13356
rect 4586 11788 4906 13300
rect 4586 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4906 11788
rect 4586 10220 4906 11732
rect 4586 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4906 10220
rect 4586 8652 4906 10164
rect 4586 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4906 8652
rect 4586 7084 4906 8596
rect 4586 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4906 7084
rect 4586 5516 4906 7028
rect 4586 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4906 5516
rect 4586 3948 4906 5460
rect 4586 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4906 3948
rect 4586 3076 4906 3892
rect 7988 15708 8308 16524
rect 7988 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8308 15708
rect 7988 14140 8308 15652
rect 7988 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8308 14140
rect 7988 12572 8308 14084
rect 7988 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8308 12572
rect 7988 11004 8308 12516
rect 7988 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8308 11004
rect 7988 9436 8308 10948
rect 7988 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8308 9436
rect 7988 7868 8308 9380
rect 7988 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8308 7868
rect 7988 6300 8308 7812
rect 7988 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8308 6300
rect 7988 4732 8308 6244
rect 7988 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8308 4732
rect 7988 3164 8308 4676
rect 7988 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8308 3164
rect 7988 3076 8308 3108
rect 11390 16492 11710 16524
rect 11390 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11710 16492
rect 11390 14924 11710 16436
rect 11390 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11710 14924
rect 11390 13356 11710 14868
rect 11390 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11710 13356
rect 11390 11788 11710 13300
rect 11390 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11710 11788
rect 11390 5516 11710 11732
rect 11390 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11710 5516
rect 11390 3948 11710 5460
rect 11390 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11710 3948
rect 11390 3076 11710 3892
rect 14792 15708 15112 16524
rect 14792 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15112 15708
rect 14792 14140 15112 15652
rect 14792 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15112 14140
rect 14792 12572 15112 14084
rect 14792 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15112 12572
rect 14792 11004 15112 12516
rect 14792 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15112 11004
rect 14792 4732 15112 10948
rect 14792 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15112 4732
rect 14792 3164 15112 4676
rect 14792 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15112 3164
rect 14792 3076 15112 3108
rect 18194 16492 18514 16524
rect 18194 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18514 16492
rect 18194 14924 18514 16436
rect 18194 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18514 14924
rect 18194 13356 18514 14868
rect 18194 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18514 13356
rect 18194 11788 18514 13300
rect 18194 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18514 11788
rect 18194 10220 18514 11732
rect 18194 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18514 10220
rect 18194 8652 18514 10164
rect 18194 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18514 8652
rect 18194 7084 18514 8596
rect 18194 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18514 7084
rect 18194 5516 18514 7028
rect 18194 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18514 5516
rect 18194 3948 18514 5460
rect 18194 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18514 3948
rect 18194 3076 18514 3892
rect 21596 15708 21916 16524
rect 21596 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21916 15708
rect 21596 14140 21916 15652
rect 21596 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21916 14140
rect 21596 12572 21916 14084
rect 21596 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21916 12572
rect 21596 11004 21916 12516
rect 21596 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21916 11004
rect 21596 9436 21916 10948
rect 21596 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21916 9436
rect 21596 7868 21916 9380
rect 21596 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21916 7868
rect 21596 6300 21916 7812
rect 21596 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21916 6300
rect 21596 4732 21916 6244
rect 21596 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21916 4732
rect 21596 3164 21916 4676
rect 21596 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21916 3164
rect 21596 3076 21916 3108
rect 24998 16492 25318 16524
rect 24998 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25318 16492
rect 24998 14924 25318 16436
rect 24998 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25318 14924
rect 24998 13356 25318 14868
rect 24998 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25318 13356
rect 24998 11788 25318 13300
rect 24998 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25318 11788
rect 24998 10220 25318 11732
rect 24998 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25318 10220
rect 24998 8652 25318 10164
rect 24998 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25318 8652
rect 24998 7084 25318 8596
rect 24998 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25318 7084
rect 24998 5516 25318 7028
rect 24998 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25318 5516
rect 24998 3948 25318 5460
rect 24998 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25318 3948
rect 24998 3076 25318 3892
rect 28400 15708 28720 16524
rect 28400 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28720 15708
rect 28400 14140 28720 15652
rect 28400 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28720 14140
rect 28400 12572 28720 14084
rect 28400 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28720 12572
rect 28400 11004 28720 12516
rect 28400 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28720 11004
rect 28400 9436 28720 10948
rect 28400 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28720 9436
rect 28400 7868 28720 9380
rect 28400 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28720 7868
rect 28400 6300 28720 7812
rect 28400 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28720 6300
rect 28400 4732 28720 6244
rect 28400 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28720 4732
rect 28400 3164 28720 4676
rect 28400 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28720 3164
rect 28400 3076 28720 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3__I
timestamp 1669390400
transform 1 0 7616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_i0_l
timestamp 1669390400
transform -1 0 10640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_i0_r
timestamp 1669390400
transform -1 0 18368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_i1_l
timestamp 1669390400
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_i1_r
timestamp 1669390400
transform 1 0 15232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_i2_l
timestamp 1669390400
transform -1 0 10192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_i2_r
timestamp 1669390400
transform 1 0 18592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_i3_l
timestamp 1669390400
transform 1 0 10416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_i3_r
timestamp 1669390400
transform 1 0 18144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_s0
timestamp 1669390400
transform 1 0 15680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_s1
timestamp 1669390400
transform 1 0 14448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_s1b
timestamp 1669390400
transform 1 0 13552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_bfg_mux_z
timestamp 1669390400
transform -1 0 14224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf_mux_I0
timestamp 1669390400
transform -1 0 7840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf_mux_I1
timestamp 1669390400
transform 1 0 3584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf_mux_I2
timestamp 1669390400
transform -1 0 3360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf_mux_I3
timestamp 1669390400
transform 1 0 7840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf_mux_S0
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf_mux_S1
timestamp 1669390400
transform 1 0 8288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 26992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform 1 0 1680 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 1904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 16912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform -1 0 24752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output7_I
timestamp 1669390400
transform 1 0 24528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3472 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55
timestamp 1669390400
transform 1 0 7504 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 8736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88
timestamp 1669390400
transform 1 0 11200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_193
timestamp 1669390400
transform 1 0 22960 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_201
timestamp 1669390400
transform 1 0 23856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_205
timestamp 1669390400
transform 1 0 24304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_229
timestamp 1669390400
transform 1 0 26992 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_237
timestamp 1669390400
transform 1 0 27888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_5
timestamp 1669390400
transform 1 0 1904 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_13
timestamp 1669390400
transform 1 0 2800 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_15
timestamp 1669390400
transform 1 0 3024 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_18
timestamp 1669390400
transform 1 0 3360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_22
timestamp 1669390400
transform 1 0 3808 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_56
timestamp 1669390400
transform 1 0 7616 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_60
timestamp 1669390400
transform 1 0 8064 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_64
timestamp 1669390400
transform 1 0 8512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_68
timestamp 1669390400
transform 1 0 8960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_231
timestamp 1669390400
transform 1 0 27216 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_239
timestamp 1669390400
transform 1 0 28112 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_69
timestamp 1669390400
transform 1 0 9072 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_72
timestamp 1669390400
transform 1 0 9408 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_104
timestamp 1669390400
transform 1 0 12992 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_107
timestamp 1669390400
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_139
timestamp 1669390400
transform 1 0 16912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_142
timestamp 1669390400
transform 1 0 17248 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_174
timestamp 1669390400
transform 1 0 20832 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_177
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_209
timestamp 1669390400
transform 1 0 24752 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_212
timestamp 1669390400
transform 1 0 25088 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_228
timestamp 1669390400
transform 1 0 26880 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_236
timestamp 1669390400
transform 1 0 27776 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_240
timestamp 1669390400
transform 1 0 28224 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_81
timestamp 1669390400
transform 1 0 10416 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_83
timestamp 1669390400
transform 1 0 10640 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_149
timestamp 1669390400
transform 1 0 18032 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_213
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_217
timestamp 1669390400
transform 1 0 25648 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_220
timestamp 1669390400
transform 1 0 25984 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_236
timestamp 1669390400
transform 1 0 27776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_240
timestamp 1669390400
transform 1 0 28224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_69
timestamp 1669390400
transform 1 0 9072 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_77
timestamp 1669390400
transform 1 0 9968 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_81
timestamp 1669390400
transform 1 0 10416 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_83
timestamp 1669390400
transform 1 0 10640 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_149
timestamp 1669390400
transform 1 0 18032 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_181
timestamp 1669390400
transform 1 0 21616 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_184
timestamp 1669390400
transform 1 0 21952 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_216
timestamp 1669390400
transform 1 0 25536 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_232
timestamp 1669390400
transform 1 0 27328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_240
timestamp 1669390400
transform 1 0 28224 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_81
timestamp 1669390400
transform 1 0 10416 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_83
timestamp 1669390400
transform 1 0 10640 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_149
timestamp 1669390400
transform 1 0 18032 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_213
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_217
timestamp 1669390400
transform 1 0 25648 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_220
timestamp 1669390400
transform 1 0 25984 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_236
timestamp 1669390400
transform 1 0 27776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_240
timestamp 1669390400
transform 1 0 28224 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_69
timestamp 1669390400
transform 1 0 9072 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_77
timestamp 1669390400
transform 1 0 9968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_83
timestamp 1669390400
transform 1 0 10640 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_149
timestamp 1669390400
transform 1 0 18032 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_152
timestamp 1669390400
transform 1 0 18368 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_168
timestamp 1669390400
transform 1 0 20160 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_180
timestamp 1669390400
transform 1 0 21504 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_184
timestamp 1669390400
transform 1 0 21952 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_200
timestamp 1669390400
transform 1 0 23744 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_208
timestamp 1669390400
transform 1 0 24640 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_225
timestamp 1669390400
transform 1 0 26544 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_229
timestamp 1669390400
transform 1 0 26992 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_237
timestamp 1669390400
transform 1 0 27888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_79
timestamp 1669390400
transform 1 0 10192 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_83
timestamp 1669390400
transform 1 0 10640 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_149
timestamp 1669390400
transform 1 0 18032 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_152
timestamp 1669390400
transform 1 0 18368 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_156
timestamp 1669390400
transform 1 0 18816 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_188
timestamp 1669390400
transform 1 0 22400 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_204
timestamp 1669390400
transform 1 0 24192 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_216
timestamp 1669390400
transform 1 0 25536 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_220
timestamp 1669390400
transform 1 0 25984 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_236
timestamp 1669390400
transform 1 0 27776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_240
timestamp 1669390400
transform 1 0 28224 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_69
timestamp 1669390400
transform 1 0 9072 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_77
timestamp 1669390400
transform 1 0 9968 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_81
timestamp 1669390400
transform 1 0 10416 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_83
timestamp 1669390400
transform 1 0 10640 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_149
timestamp 1669390400
transform 1 0 18032 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_181
timestamp 1669390400
transform 1 0 21616 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_184
timestamp 1669390400
transform 1 0 21952 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_216
timestamp 1669390400
transform 1 0 25536 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_232
timestamp 1669390400
transform 1 0 27328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_240
timestamp 1669390400
transform 1 0 28224 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_81
timestamp 1669390400
transform 1 0 10416 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_83
timestamp 1669390400
transform 1 0 10640 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_149
timestamp 1669390400
transform 1 0 18032 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_213
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_217
timestamp 1669390400
transform 1 0 25648 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_220
timestamp 1669390400
transform 1 0 25984 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_236
timestamp 1669390400
transform 1 0 27776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_240
timestamp 1669390400
transform 1 0 28224 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_69
timestamp 1669390400
transform 1 0 9072 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_72
timestamp 1669390400
transform 1 0 9408 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_88
timestamp 1669390400
transform 1 0 11200 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_96
timestamp 1669390400
transform 1 0 12096 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_100
timestamp 1669390400
transform 1 0 12544 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_104
timestamp 1669390400
transform 1 0 12992 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_107
timestamp 1669390400
transform 1 0 13328 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_111
timestamp 1669390400
transform 1 0 13776 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_115
timestamp 1669390400
transform 1 0 14224 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_119
timestamp 1669390400
transform 1 0 14672 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_123
timestamp 1669390400
transform 1 0 15120 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_126
timestamp 1669390400
transform 1 0 15456 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_130
timestamp 1669390400
transform 1 0 15904 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_138
timestamp 1669390400
transform 1 0 16800 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_142
timestamp 1669390400
transform 1 0 17248 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_174
timestamp 1669390400
transform 1 0 20832 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_177
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_209
timestamp 1669390400
transform 1 0 24752 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_212
timestamp 1669390400
transform 1 0 25088 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_228
timestamp 1669390400
transform 1 0 26880 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_236
timestamp 1669390400
transform 1 0 27776 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_240
timestamp 1669390400
transform 1 0 28224 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_5
timestamp 1669390400
transform 1 0 1904 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_69
timestamp 1669390400
transform 1 0 9072 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_231
timestamp 1669390400
transform 1 0 27216 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_239
timestamp 1669390400
transform 1 0 28112 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_19
timestamp 1669390400
transform 1 0 3472 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_45
timestamp 1669390400
transform 1 0 6384 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_49
timestamp 1669390400
transform 1 0 6832 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_54
timestamp 1669390400
transform 1 0 7392 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_58
timestamp 1669390400
transform 1 0 7840 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_90
timestamp 1669390400
transform 1 0 11424 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_211
timestamp 1669390400
transform 1 0 24976 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_227
timestamp 1669390400
transform 1 0 26768 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_235
timestamp 1669390400
transform 1 0 27664 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_239
timestamp 1669390400
transform 1 0 28112 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_105
timestamp 1669390400
transform 1 0 13104 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_121
timestamp 1669390400
transform 1 0 14896 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_129
timestamp 1669390400
transform 1 0 15792 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_133
timestamp 1669390400
transform 1 0 16240 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_138
timestamp 1669390400
transform 1 0 16800 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_147
timestamp 1669390400
transform 1 0 17808 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_211
timestamp 1669390400
transform 1 0 24976 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_231
timestamp 1669390400
transform 1 0 27216 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_239
timestamp 1669390400
transform 1 0 28112 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1669390400
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_211
timestamp 1669390400
transform 1 0 24976 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_227
timestamp 1669390400
transform 1 0 26768 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_235
timestamp 1669390400
transform 1 0 27664 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_239
timestamp 1669390400
transform 1 0 28112 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_231
timestamp 1669390400
transform 1 0 27216 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_239
timestamp 1669390400
transform 1 0 28112 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_18
timestamp 1669390400
transform 1 0 3360 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_26
timestamp 1669390400
transform 1 0 4256 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_30
timestamp 1669390400
transform 1 0 4704 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_54
timestamp 1669390400
transform 1 0 7392 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_72
timestamp 1669390400
transform 1 0 9408 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_104
timestamp 1669390400
transform 1 0 12992 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_107
timestamp 1669390400
transform 1 0 13328 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_123
timestamp 1669390400
transform 1 0 15120 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_131
timestamp 1669390400
transform 1 0 16016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_135
timestamp 1669390400
transform 1 0 16464 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_139
timestamp 1669390400
transform 1 0 16912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_142
timestamp 1669390400
transform 1 0 17248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_144
timestamp 1669390400
transform 1 0 17472 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_170
timestamp 1669390400
transform 1 0 20384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_174
timestamp 1669390400
transform 1 0 20832 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_177
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_193
timestamp 1669390400
transform 1 0 22960 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_201
timestamp 1669390400
transform 1 0 23856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_205
timestamp 1669390400
transform 1 0 24304 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_209
timestamp 1669390400
transform 1 0 24752 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_212
timestamp 1669390400
transform 1 0 25088 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_227
timestamp 1669390400
transform 1 0 26768 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_235
timestamp 1669390400
transform 1 0 27664 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_239
timestamp 1669390400
transform 1 0 28112 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 28560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 10976 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 17808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 28560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 10976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 17808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 10976 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 17808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 28560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 10976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 17808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 10976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 17808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 28560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 10976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 17808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 10976 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 17808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 28560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 28560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_52
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_53
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_54
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_55
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_56
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_57
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_58
timestamp 1669390400
transform 1 0 9184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_59
timestamp 1669390400
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_60
timestamp 1669390400
transform 1 0 17024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_61
timestamp 1669390400
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_62
timestamp 1669390400
transform 1 0 24864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_63
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_64
timestamp 1669390400
transform 1 0 25760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_65
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_66
timestamp 1669390400
transform 1 0 21728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_67
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_68
timestamp 1669390400
transform 1 0 25760 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_69
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_70
timestamp 1669390400
transform 1 0 21728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_71
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_72
timestamp 1669390400
transform 1 0 25760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_73
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_74
timestamp 1669390400
transform 1 0 21728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_75
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_76
timestamp 1669390400
transform 1 0 25760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_77
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_78
timestamp 1669390400
transform 1 0 9184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_79
timestamp 1669390400
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_80
timestamp 1669390400
transform 1 0 17024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_81
timestamp 1669390400
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_82
timestamp 1669390400
transform 1 0 24864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_83
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_84
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_85
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1669390400
transform 1 0 9184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1669390400
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1669390400
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1669390400
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1669390400
transform 1 0 24864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 16800 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3_
timestamp 1669390400
transform 1 0 6944 0 1 12544
box -86 -86 534 870
use gf180mcu_mux  bfg_mux
timestamp 0
transform 1 0 13090 0 1 8062
box 0 -49 2478 709
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  gf_mux dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7616 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 26544 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 1680 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform 1 0 1680 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform 1 0 5600 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input5 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 20384 0 1 15680
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input6
timestamp 1669390400
transform -1 0 26992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output7 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 25200 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output8
timestamp 1669390400
transform 1 0 11424 0 1 3136
box -86 -86 1654 870
<< labels >>
flabel metal2 s 29568 19200 29680 19800 0 FreeSans 448 90 0 0 bfg_out
port 0 nsew signal tristate
flabel metal2 s 12096 200 12208 800 0 FreeSans 448 90 0 0 gf_out
port 1 nsew signal tristate
flabel metal3 s 29200 7392 29800 7504 0 FreeSans 448 0 0 0 i0
port 2 nsew signal input
flabel metal3 s 200 12096 800 12208 0 FreeSans 448 0 0 0 i1
port 3 nsew signal input
flabel metal2 s 0 200 112 800 0 FreeSans 448 90 0 0 i2
port 4 nsew signal input
flabel metal2 s 4704 19200 4816 19800 0 FreeSans 448 90 0 0 i3
port 5 nsew signal input
flabel metal2 s 17472 19200 17584 19800 0 FreeSans 448 90 0 0 s0
port 6 nsew signal input
flabel metal2 s 24864 200 24976 800 0 FreeSans 448 90 0 0 s1
port 7 nsew signal input
flabel metal4 s 4586 3076 4906 16524 0 FreeSans 1280 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 11390 3076 11710 16524 0 FreeSans 1280 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 18194 3076 18514 16524 0 FreeSans 1280 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 24998 3076 25318 16524 0 FreeSans 1280 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 7988 3076 8308 16524 0 FreeSans 1280 90 0 0 vss
port 9 nsew ground bidirectional
flabel metal4 s 14792 3076 15112 16524 0 FreeSans 1280 90 0 0 vss
port 9 nsew ground bidirectional
flabel metal4 s 21596 3076 21916 16524 0 FreeSans 1280 90 0 0 vss
port 9 nsew ground bidirectional
flabel metal4 s 28400 3076 28720 16524 0 FreeSans 1280 90 0 0 vss
port 9 nsew ground bidirectional
rlabel metal1 23184 10192 23184 10192 0 vdd
rlabel metal1 23264 9408 23264 9408 0 vss
rlabel metal1 13888 8826 13888 8826 0 _0_
rlabel metal2 13608 12096 13608 12096 0 _1_
rlabel metal2 26488 16968 26488 16968 0 bfg_out
rlabel metal2 12152 2198 12152 2198 0 gf_out
rlabel metal2 26936 7728 26936 7728 0 i0
rlabel metal3 1246 12152 1246 12152 0 i1
rlabel metal2 1960 2968 1960 2968 0 i2
rlabel metal2 4984 16632 4984 16632 0 i3
rlabel metal2 4424 4368 4424 4368 0 net1
rlabel metal3 4424 4312 4424 4312 0 net2
rlabel metal2 7448 5656 7448 5656 0 net3
rlabel metal2 7896 4704 7896 4704 0 net4
rlabel metal2 7112 4256 7112 4256 0 net5
rlabel metal3 7168 4312 7168 4312 0 net6
rlabel metal2 24584 15680 24584 15680 0 net7
rlabel metal2 6440 3976 6440 3976 0 net8
rlabel metal3 17192 16184 17192 16184 0 s0
rlabel metal2 24808 3416 24808 3416 0 s1
<< properties >>
string FIXED_BBOX 0 0 30000 20000
<< end >>
